VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
   DATABASE MICRONS 1000 ;
END UNITS

MACRO h3
   CLASS BLOCK ;
   FOREIGN h3 ;
   ORIGIN 0 0 ;
   SIZE 549.2 BY 296 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1005_n_65753
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 76.55 0.51 76.65 ;
      END
   END FE_OFN1005_n_65753

   PIN FE_OFN1022_n_3701
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.35 0.51 29.45 ;
      END
   END FE_OFN1022_n_3701

   PIN FE_OFN1051_n_5643
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 243.75 0.51 243.85 ;
      END
   END FE_OFN1051_n_5643

   PIN FE_OFN106_n_95123
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.95 0.51 112.05 ;
      END
   END FE_OFN106_n_95123

   PIN FE_OFN1075_n_116
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 23.6 0 23.8 0.255 ;
      END
   END FE_OFN1075_n_116

   PIN FE_OFN1095_g303299_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.55 0.51 16.65 ;
      END
   END FE_OFN1095_g303299_p

   PIN FE_OFN1121_n_4882
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 243.95 0.51 244.05 ;
      END
   END FE_OFN1121_n_4882

   PIN FE_OFN1203_n_118585
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 178.2 0 178.4 0.255 ;
      END
   END FE_OFN1203_n_118585

   PIN FE_OFN1215_n_3935
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.75 0.51 16.85 ;
      END
   END FE_OFN1215_n_3935

   PIN FE_OFN1225_n_6583
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.65 0 83.75 0.51 ;
      END
   END FE_OFN1225_n_6583

   PIN FE_OFN1228_n_3045
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.25 0 14.35 0.51 ;
      END
   END FE_OFN1228_n_3045

   PIN FE_OFN1431_n_22026
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 40.45 0 40.55 0.51 ;
      END
   END FE_OFN1431_n_22026

   PIN FE_OFN1534_n_4068
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.95 0.51 17.05 ;
      END
   END FE_OFN1534_n_4068

   PIN FE_OFN1551_n_13938
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.95 0.51 33.05 ;
      END
   END FE_OFN1551_n_13938

   PIN FE_OFN1579_n_3047
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.15 0.51 17.25 ;
      END
   END FE_OFN1579_n_3047

   PIN FE_OFN1625_n_3863
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.35 0.51 17.45 ;
      END
   END FE_OFN1625_n_3863

   PIN FE_OFN1667_n_66371
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.85 0 86.95 0.51 ;
      END
   END FE_OFN1667_n_66371

   PIN FE_OFN1863_n_4923
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.55 0.51 17.65 ;
      END
   END FE_OFN1863_n_4923

   PIN FE_OFN1930_n_18862
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.75 0.51 17.85 ;
      END
   END FE_OFN1930_n_18862

   PIN FE_OFN1959_n_6873
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 94.45 0 94.55 0.51 ;
      END
   END FE_OFN1959_n_6873

   PIN FE_OFN2010_n_27918
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.85 0 57.95 0.51 ;
      END
   END FE_OFN2010_n_27918

   PIN FE_OFN2014_n_23906
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 195.75 0.51 195.85 ;
      END
   END FE_OFN2014_n_23906

   PIN FE_OFN2148_n_118596
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.95 0.51 13.05 ;
      END
   END FE_OFN2148_n_118596

   PIN FE_OFN2171_n_117298
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 165.85 0 165.95 0.51 ;
      END
   END FE_OFN2171_n_117298

   PIN FE_OFN2175_n_21905
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 12.95 0.51 13.05 ;
      END
   END FE_OFN2175_n_21905

   PIN FE_OFN2254_n_23876
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 13.15 0.51 13.25 ;
      END
   END FE_OFN2254_n_23876

   PIN FE_OFN2334_n_23919
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 11.35 0.51 11.45 ;
      END
   END FE_OFN2334_n_23919

   PIN FE_OFN2352_n_27890
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 103.65 0 103.75 0.51 ;
      END
   END FE_OFN2352_n_27890

   PIN FE_OFN2353_n_19056
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 17.95 0.51 18.05 ;
      END
   END FE_OFN2353_n_19056

   PIN FE_OFN2395_n_61534
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.15 0.51 18.25 ;
      END
   END FE_OFN2395_n_61534

   PIN FE_OFN2397_n_4104
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.75 0.51 23.85 ;
      END
   END FE_OFN2397_n_4104

   PIN FE_OFN2400_n_18228
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 22.95 0.51 23.05 ;
      END
   END FE_OFN2400_n_18228

   PIN FE_OFN2418_n_26365
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 52.85 0 52.95 0.51 ;
      END
   END FE_OFN2418_n_26365

   PIN FE_OFN2419_n_25888
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 172.35 0.51 172.45 ;
      END
   END FE_OFN2419_n_25888

   PIN FE_OFN2473_n_117820
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 330.45 0 330.55 0.51 ;
      END
   END FE_OFN2473_n_117820

   PIN FE_OFN2484_n_25794
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 13.35 0.51 13.45 ;
      END
   END FE_OFN2484_n_25794

   PIN FE_OFN2502_n_5437
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 79.05 0 79.15 0.51 ;
      END
   END FE_OFN2502_n_5437

   PIN FE_OFN2505_n_4918
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 195.95 0.51 196.05 ;
      END
   END FE_OFN2505_n_4918

   PIN FE_OFN2678_n_23958
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 255.75 0.51 255.85 ;
      END
   END FE_OFN2678_n_23958

   PIN FE_OFN2701_n_2549
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 51.15 0.51 51.25 ;
      END
   END FE_OFN2701_n_2549

   PIN FE_OFN2720_n_25980
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.15 0.51 112.25 ;
      END
   END FE_OFN2720_n_25980

   PIN FE_OFN2787_n_5684
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.35 0.51 112.45 ;
      END
   END FE_OFN2787_n_5684

   PIN FE_OFN2790_n_4079
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 5.25 0 5.35 0.51 ;
      END
   END FE_OFN2790_n_4079

   PIN FE_OFN287_n_76853
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.65 0 24.75 0.51 ;
      END
   END FE_OFN287_n_76853

   PIN FE_OFN2929_n_4064
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 26.05 0 26.15 0.51 ;
      END
   END FE_OFN2929_n_4064

   PIN FE_OFN2976_n_65768
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.15 0.51 111.25 ;
      END
   END FE_OFN2976_n_65768

   PIN FE_OFN3004_n_4088
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 12.65 0 12.75 0.51 ;
      END
   END FE_OFN3004_n_4088

   PIN FE_OFN3018_n_69766
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 306.25 0 306.35 0.51 ;
      END
   END FE_OFN3018_n_69766

   PIN FE_OFN3050_n_3016
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.15 0.51 63.25 ;
      END
   END FE_OFN3050_n_3016

   PIN FE_OFN3096_n_4811
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.55 0.51 25.65 ;
      END
   END FE_OFN3096_n_4811

   PIN FE_OFN3163_n_2780
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 2.25 0 2.35 0.51 ;
      END
   END FE_OFN3163_n_2780

   PIN FE_OFN3206_n_32181
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 172.25 0 172.35 0.51 ;
      END
   END FE_OFN3206_n_32181

   PIN FE_OFN3230_n_3189
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.45 0 5.55 0.51 ;
      END
   END FE_OFN3230_n_3189

   PIN FE_OFN3235_n_2155
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.45 0 10.55 0.51 ;
      END
   END FE_OFN3235_n_2155

   PIN FE_OFN3241_n_4790
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.75 0.51 25.85 ;
      END
   END FE_OFN3241_n_4790

   PIN FE_OFN325_n_70684
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 294.85 0 294.95 0.51 ;
      END
   END FE_OFN325_n_70684

   PIN FE_OFN327_n_70685
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.65 0 318.75 0.51 ;
      END
   END FE_OFN327_n_70685

   PIN FE_OFN3364_n_25895
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 208.35 0.51 208.45 ;
      END
   END FE_OFN3364_n_25895

   PIN FE_OFN3366_n_5443
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 255.95 0.51 256.05 ;
      END
   END FE_OFN3366_n_5443

   PIN FE_OFN3464_n_67106
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.65 295.49 127.75 296 ;
      END
   END FE_OFN3464_n_67106

   PIN FE_OFN3486_n_1596
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 13.55 0.51 13.65 ;
      END
   END FE_OFN3486_n_1596

   PIN FE_OFN3517_n_23820
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 33.15 0.51 33.25 ;
      END
   END FE_OFN3517_n_23820

   PIN FE_OFN3531_n_19107
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.7 0.255 24.9 ;
      END
   END FE_OFN3531_n_19107

   PIN FE_OFN3549_n_7898
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 33.35 0.51 33.45 ;
      END
   END FE_OFN3549_n_7898

   PIN FE_OFN3617_n_18380
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 13.75 0.51 13.85 ;
      END
   END FE_OFN3617_n_18380

   PIN FE_OFN3628_n_4557
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.55 0.51 88.65 ;
      END
   END FE_OFN3628_n_4557

   PIN FE_OFN3720_n_4799
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 11.55 0.51 11.65 ;
      END
   END FE_OFN3720_n_4799

   PIN FE_OFN3800_n_23840
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.35 0.51 18.45 ;
      END
   END FE_OFN3800_n_23840

   PIN FE_OFN3910_n_5532
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 244.15 0.51 244.25 ;
      END
   END FE_OFN3910_n_5532

   PIN FE_OFN4090_n_2663
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 18.15 0.51 18.25 ;
      END
   END FE_OFN4090_n_2663

   PIN FE_OFN4798_n_21953
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.55 0.51 18.65 ;
      END
   END FE_OFN4798_n_21953

   PIN FE_OFN666_n_31829
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 160.65 0 160.75 0.51 ;
      END
   END FE_OFN666_n_31829

   PIN FE_OFN693_n_27625
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.65 0 34.75 0.51 ;
      END
   END FE_OFN693_n_27625

   PIN FE_OFN715_n_24030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 13.45 0 13.55 0.51 ;
      END
   END FE_OFN715_n_24030

   PIN FE_OFN737_n_4131
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.75 0.51 18.85 ;
      END
   END FE_OFN737_n_4131

   PIN FE_OFN847_n_4294
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 18.95 0.51 19.05 ;
      END
   END FE_OFN847_n_4294

   PIN FE_OFN848_n_4958
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 51.35 0.51 51.45 ;
      END
   END FE_OFN848_n_4958

   PIN FE_OFN853_n_3353
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 19.15 0.51 19.25 ;
      END
   END FE_OFN853_n_3353

   PIN FE_OFN911_n_21872
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 18.35 0.51 18.45 ;
      END
   END FE_OFN911_n_21872

   PIN FE_OFN948_n_3795
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.95 0.51 26.05 ;
      END
   END FE_OFN948_n_3795

   PIN FE_OFN965_n_25771
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 19.35 0.51 19.45 ;
      END
   END FE_OFN965_n_25771

   PIN FE_OFN973_n_63299
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 19.55 0.51 19.65 ;
      END
   END FE_OFN973_n_63299

   PIN FE_OFN975_n_2435
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.95 0.51 24.05 ;
      END
   END FE_OFN975_n_2435

   PIN g205805_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.05 0 232.15 0.51 ;
      END
   END g205805_da

   PIN g221053_u1_o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.05 295.49 56.15 296 ;
      END
   END g221053_u1_o

   PIN g222840_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 33.55 0.51 33.65 ;
      END
   END g222840_p

   PIN g229165_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.25 0 320.35 0.51 ;
      END
   END g229165_p

   PIN g229250_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.45 0 320.55 0.51 ;
      END
   END g229250_p

   PIN g229781_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 73.25 0 73.35 0.51 ;
      END
   END g229781_p

   PIN g231281_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.35 0.51 63.45 ;
      END
   END g231281_p

   PIN g233246_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.05 0 36.15 0.51 ;
      END
   END g233246_p

   PIN g233290_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.75 0.51 51.85 ;
      END
   END g233290_p

   PIN g233318_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.85 0 78.95 0.51 ;
      END
   END g233318_p

   PIN g233379_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 75.05 0 75.15 0.51 ;
      END
   END g233379_p

   PIN g233525_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.55 0.51 124.65 ;
      END
   END g233525_p

   PIN g233666_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.35 0.51 39.45 ;
      END
   END g233666_p

   PIN g233787_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.55 0.51 28.65 ;
      END
   END g233787_p

   PIN g235027_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 61.65 0 61.75 0.51 ;
      END
   END g235027_p

   PIN g235236_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 66.45 0 66.55 0.51 ;
      END
   END g235236_p

   PIN g235278_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 62.25 0 62.35 0.51 ;
      END
   END g235278_p

   PIN g235292_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.25 0 78.35 0.51 ;
      END
   END g235292_p

   PIN g235499_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 172.55 0.51 172.65 ;
      END
   END g235499_p

   PIN g235503_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 61.05 0 61.15 0.51 ;
      END
   END g235503_p

   PIN g236596_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35.05 0 35.15 0.51 ;
      END
   END g236596_da

   PIN g236596_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.25 0 29.35 0.51 ;
      END
   END g236596_db

   PIN g264946_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.05 0 271.15 0.51 ;
      END
   END g264946_da

   PIN g264946_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.85 0 271.95 0.51 ;
      END
   END g264946_db

   PIN g265666_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.65 0 292.75 0.51 ;
      END
   END g265666_p

   PIN g265686_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 295.25 0 295.35 0.51 ;
      END
   END g265686_p

   PIN g265687_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.45 0 294.55 0.51 ;
      END
   END g265687_p

   PIN g266335_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.45 0 271.55 0.51 ;
      END
   END g266335_p

   PIN g267264_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 192.45 0 192.55 0.51 ;
      END
   END g267264_da

   PIN g267734_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 207.85 0 207.95 0.51 ;
      END
   END g267734_p

   PIN g267768_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 204.25 0 204.35 0.51 ;
      END
   END g267768_p

   PIN g267963_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 202.05 0 202.15 0.51 ;
      END
   END g267963_p

   PIN g269325_p1
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 332.05 0 332.15 0.51 ;
      END
   END g269325_p1

   PIN g270287_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 212.45 0 212.55 0.51 ;
      END
   END g270287_p

   PIN g270719_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 132.65 0 132.75 0.51 ;
      END
   END g270719_p

   PIN g270759_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 193.25 0 193.35 0.51 ;
      END
   END g270759_da

   PIN g270759_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 193.25 0 193.35 0.51 ;
      END
   END g270759_db

   PIN g271925_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 94.25 0 94.35 0.51 ;
      END
   END g271925_p

   PIN g271962_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.65 0 100.75 0.51 ;
      END
   END g271962_p

   PIN g271983_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 95.65 0 95.75 0.51 ;
      END
   END g271983_p

   PIN g272146_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.05 0 103.15 0.51 ;
      END
   END g272146_p

   PIN g273791_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.55 0.51 63.65 ;
      END
   END g273791_p

   PIN g274959_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 46.85 0 46.95 0.51 ;
      END
   END g274959_p

   PIN g275109_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 24.85 0 24.95 0.51 ;
      END
   END g275109_sb

   PIN g275315_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.85 295.49 28.95 296 ;
      END
   END g275315_da

   PIN g275315_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 32.25 295.49 32.35 296 ;
      END
   END g275315_db

   PIN g279718_p2
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 220.35 0.51 220.45 ;
      END
   END g279718_p2

   PIN g279854_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 196.15 0.51 196.25 ;
      END
   END g279854_p

   PIN g280604_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 184.55 0.51 184.65 ;
      END
   END g280604_p

   PIN g281129_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.85 0 11.95 0.51 ;
      END
   END g281129_p

   PIN g302688_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.65 0 5.75 0.51 ;
      END
   END g302688_p

   PIN g302697_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 17.65 0 17.75 0.51 ;
      END
   END g302697_p

   PIN g302698_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 11.75 0.51 11.85 ;
      END
   END g302698_p

   PIN g302705_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.65 0 26.75 0.51 ;
      END
   END g302705_p

   PIN g303296_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 10.95 0.51 11.05 ;
      END
   END g303296_p

   PIN g303330_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.55 0.51 29.65 ;
      END
   END g303330_p

   PIN g303332_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 42.25 0 42.35 0.51 ;
      END
   END g303332_p

   PIN g303358_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 11.95 0.51 12.05 ;
      END
   END g303358_p

   PIN g304265_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.85 0 8.95 0.51 ;
      END
   END g304265_p

   PIN g304267_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.25 0 28.35 0.51 ;
      END
   END g304267_p

   PIN g304295_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 13.25 0 13.35 0.51 ;
      END
   END g304295_p

   PIN g304307_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.75 0.51 63.85 ;
      END
   END g304307_p

   PIN g304312_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.05 0 7.15 0.51 ;
      END
   END g304312_p

   PIN g304735_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 38.95 0.51 39.05 ;
      END
   END g304735_p

   PIN g304777_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.75 0.51 29.85 ;
      END
   END g304777_p

   PIN g322260_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.85 0 211.95 0.51 ;
      END
   END g322260_p

   PIN g322487_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.25 0 320.35 0.51 ;
      END
   END g322487_p

   PIN g322619_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.85 0 159.95 0.51 ;
      END
   END g322619_da

   PIN g322619_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 235.65 0 235.75 0.51 ;
      END
   END g322619_db

   PIN n_1057
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 19.75 0.51 19.85 ;
      END
   END n_1057

   PIN n_108861
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.75 0.51 124.85 ;
      END
   END n_108861

   PIN n_109000
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 19.95 0.51 20.05 ;
      END
   END n_109000

   PIN n_109172
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.25 0 2.35 0.51 ;
      END
   END n_109172

   PIN n_109184
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 81.65 0 81.75 0.51 ;
      END
   END n_109184

   PIN n_1098
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.15 0.51 52.25 ;
      END
   END n_1098

   PIN n_112975
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 372.45 0 372.55 0.51 ;
      END
   END n_112975

   PIN n_112976
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 367.85 0 367.95 0.51 ;
      END
   END n_112976

   PIN n_113031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 227.05 0 227.15 0.51 ;
      END
   END n_113031

   PIN n_116915
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.85 0 55.95 0.51 ;
      END
   END n_116915

   PIN n_116916
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 26.6 0 26.8 0.255 ;
      END
   END n_116916

   PIN n_116953
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 52.25 0 52.35 0.51 ;
      END
   END n_116953

   PIN n_117338
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 25.15 0.51 25.25 ;
      END
   END n_117338

   PIN n_117342
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 18.55 0.51 18.65 ;
      END
   END n_117342

   PIN n_117601
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 235.05 0 235.15 0.51 ;
      END
   END n_117601

   PIN n_117819
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 332.65 0 332.75 0.51 ;
      END
   END n_117819

   PIN n_118320
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 115.45 0 115.55 0.51 ;
      END
   END n_118320

   PIN n_118334
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.85 0 163.95 0.51 ;
      END
   END n_118334

   PIN n_118459
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 43.45 0 43.55 0.51 ;
      END
   END n_118459

   PIN n_118597
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.85 295.49 17.95 296 ;
      END
   END n_118597

   PIN n_118744
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 184.75 0.51 184.85 ;
      END
   END n_118744

   PIN n_118754
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 186.65 0 186.75 0.51 ;
      END
   END n_118754

   PIN n_126138
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.95 0.51 52.05 ;
      END
   END n_126138

   PIN n_1264
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.25 0 7.35 0.51 ;
      END
   END n_1264

   PIN n_1278
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.65 0 11.75 0.51 ;
      END
   END n_1278

   PIN n_13895
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 16.65 0 16.75 0.51 ;
      END
   END n_13895

   PIN n_140823
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 194.25 0 194.35 0.51 ;
      END
   END n_140823

   PIN n_1464
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.25 0 15.35 0.51 ;
      END
   END n_1464

   PIN n_1469
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.45 0 2.55 0.51 ;
      END
   END n_1469

   PIN n_1482
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 5.05 0 5.15 0.51 ;
      END
   END n_1482

   PIN n_1507
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 18.75 0.51 18.85 ;
      END
   END n_1507

   PIN n_1511
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.65 0 6.75 0.51 ;
      END
   END n_1511

   PIN n_151614
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 1.05 0 1.15 0.51 ;
      END
   END n_151614

   PIN n_1599
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.95 0.51 63.05 ;
      END
   END n_1599

   PIN n_162433
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 196.35 0.51 196.45 ;
      END
   END n_162433

   PIN n_1790
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 39.15 0.51 39.25 ;
      END
   END n_1790

   PIN n_18375
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 207.55 0.51 207.65 ;
      END
   END n_18375

   PIN n_183956
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 58.25 0 58.35 0.51 ;
      END
   END n_183956

   PIN n_1867
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 21.95 0.51 22.05 ;
      END
   END n_1867

   PIN n_1932
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.05 0 6.15 0.51 ;
      END
   END n_1932

   PIN n_1952
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.35 0.51 34.45 ;
      END
   END n_1952

   PIN n_19942
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 208.55 0.51 208.65 ;
      END
   END n_19942

   PIN n_19943
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 207.75 0.51 207.85 ;
      END
   END n_19943

   PIN n_19987
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 13.35 0.51 13.45 ;
      END
   END n_19987

   PIN n_20051
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 11.15 0.51 11.25 ;
      END
   END n_20051

   PIN n_2049
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.85 0 14.95 0.51 ;
      END
   END n_2049

   PIN n_20823
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 13.05 0 13.15 0.51 ;
      END
   END n_20823

   PIN n_20967
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 196.55 0.51 196.65 ;
      END
   END n_20967

   PIN n_21560
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.05 0 4.15 0.51 ;
      END
   END n_21560

   PIN n_21836
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 19.45 0 19.55 0.51 ;
      END
   END n_21836

   PIN n_21898
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 63.15 0.51 63.25 ;
      END
   END n_21898

   PIN n_21970
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.85 0 19.95 0.51 ;
      END
   END n_21970

   PIN n_21978
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.05 0 56.15 0.51 ;
      END
   END n_21978

   PIN n_21997
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.65 0 2.75 0.51 ;
      END
   END n_21997

   PIN n_22074
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.35 0.51 36.45 ;
      END
   END n_22074

   PIN n_22077
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.85 0 16.95 0.51 ;
      END
   END n_22077

   PIN n_22109
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.25 0 23.35 0.51 ;
      END
   END n_22109

   PIN n_22116
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 54.65 0 54.75 0.51 ;
      END
   END n_22116

   PIN n_22254
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.35 0.51 32.45 ;
      END
   END n_22254

   PIN n_22267
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.05 0 26.15 0.51 ;
      END
   END n_22267

   PIN n_22272
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.05 0 2.15 0.51 ;
      END
   END n_22272

   PIN n_22339
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.25 0 26.35 0.51 ;
      END
   END n_22339

   PIN n_22384
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 17.2 0 17.4 0.255 ;
      END
   END n_22384

   PIN n_22477
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.55 0.51 33.65 ;
      END
   END n_22477

   PIN n_22600
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 54.85 0 54.95 0.51 ;
      END
   END n_22600

   PIN n_22668
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 39.35 0.51 39.45 ;
      END
   END n_22668

   PIN n_22760
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.05 0 17.15 0.51 ;
      END
   END n_22760

   PIN n_22793
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.45 0 17.55 0.51 ;
      END
   END n_22793

   PIN n_22810
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.65 0 17.75 0.51 ;
      END
   END n_22810

   PIN n_22832
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 51.55 0.51 51.65 ;
      END
   END n_22832

   PIN n_22938
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.65 0 20.75 0.51 ;
      END
   END n_22938

   PIN n_23072
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.85 0 15.95 0.51 ;
      END
   END n_23072

   PIN n_23082
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 21.35 0.51 21.45 ;
      END
   END n_23082

   PIN n_23089
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.55 0.51 31.65 ;
      END
   END n_23089

   PIN n_23126
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 16.85 0 16.95 0.51 ;
      END
   END n_23126

   PIN n_23209
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 13.05 0 13.15 0.51 ;
      END
   END n_23209

   PIN n_23215
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.55 0.51 36.65 ;
      END
   END n_23215

   PIN n_2327
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.45 0 21.55 0.51 ;
      END
   END n_2327

   PIN n_23391
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 19.05 0 19.15 0.51 ;
      END
   END n_23391

   PIN n_23480
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.45 0 20.55 0.51 ;
      END
   END n_23480

   PIN n_23488
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 20.55 0.51 20.65 ;
      END
   END n_23488

   PIN n_23559
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 26.95 0.51 27.05 ;
      END
   END n_23559

   PIN n_23605
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.45 0 19.55 0.51 ;
      END
   END n_23605

   PIN n_23607
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.25 0 21.35 0.51 ;
      END
   END n_23607

   PIN n_23658
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.05 0 23.15 0.51 ;
      END
   END n_23658

   PIN n_23760
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 76.75 0.51 76.85 ;
      END
   END n_23760

   PIN n_23795
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.15 0.51 26.25 ;
      END
   END n_23795

   PIN n_23805
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 63.35 0.51 63.45 ;
      END
   END n_23805

   PIN n_23889
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 404.05 295.49 404.15 296 ;
      END
   END n_23889

   PIN n_23929
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 524.05 0 524.15 0.51 ;
      END
   END n_23929

   PIN n_24160
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 33.75 0.51 33.85 ;
      END
   END n_24160

   PIN n_24271
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 75.95 0.51 76.05 ;
      END
   END n_24271

   PIN n_24308
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.65 0 3.75 0.51 ;
      END
   END n_24308

   PIN n_24929
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.7 0.255 22.9 ;
      END
   END n_24929

   PIN n_25559
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.75 0.51 28.85 ;
      END
   END n_25559

   PIN n_25809
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 256.15 0.51 256.25 ;
      END
   END n_25809

   PIN n_25811
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.55 0.51 112.65 ;
      END
   END n_25811

   PIN n_25812
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 171.75 0.51 171.85 ;
      END
   END n_25812

   PIN n_25904
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.55 0.51 9.65 ;
      END
   END n_25904

   PIN n_25932
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.45 0 174.55 0.51 ;
      END
   END n_25932

   PIN n_25934
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 256.35 0.51 256.45 ;
      END
   END n_25934

   PIN n_25939
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 244.35 0.51 244.45 ;
      END
   END n_25939

   PIN n_25994
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 76.95 0.51 77.05 ;
      END
   END n_25994

   PIN n_26053
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 279.95 0.51 280.05 ;
      END
   END n_26053

   PIN n_26162
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.65 0 12.75 0.51 ;
      END
   END n_26162

   PIN n_26171
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.9 0.255 47.1 ;
      END
   END n_26171

   PIN n_26172
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.75 0.51 43.85 ;
      END
   END n_26172

   PIN n_26188
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 256.55 0.51 256.65 ;
      END
   END n_26188

   PIN n_26255
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.75 0.51 44.85 ;
      END
   END n_26255

   PIN n_26333
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 7.65 0 7.75 0.51 ;
      END
   END n_26333

   PIN n_26360
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.35 0.51 9.45 ;
      END
   END n_26360

   PIN n_26362
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.95 0.51 64.05 ;
      END
   END n_26362

   PIN n_26373
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 47.35 0.51 47.45 ;
      END
   END n_26373

   PIN n_26495
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.35 0.51 45.45 ;
      END
   END n_26495

   PIN n_26507
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.95 0.51 10.05 ;
      END
   END n_26507

   PIN n_26533
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.15 0.51 44.25 ;
      END
   END n_26533

   PIN n_26619
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 25.55 0.51 25.65 ;
      END
   END n_26619

   PIN n_26627
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.15 0.51 50.25 ;
      END
   END n_26627

   PIN n_26634
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 100.15 0.51 100.25 ;
      END
   END n_26634

   PIN n_26662
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 47.55 0.51 47.65 ;
      END
   END n_26662

   PIN n_26750
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.15 0.51 64.25 ;
      END
   END n_26750

   PIN n_26760
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.55 0.51 45.65 ;
      END
   END n_26760

   PIN n_26773
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.75 0.51 62.85 ;
      END
   END n_26773

   PIN n_26775
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 41.55 0.51 41.65 ;
      END
   END n_26775

   PIN n_26929
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 21.75 0.51 21.85 ;
      END
   END n_26929

   PIN n_27125
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 78.05 0 78.15 0.51 ;
      END
   END n_27125

   PIN n_27252
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 25.75 0.51 25.85 ;
      END
   END n_27252

   PIN n_27259
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.75 0.51 45.85 ;
      END
   END n_27259

   PIN n_27388
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 36.95 0.51 37.05 ;
      END
   END n_27388

   PIN n_27391
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 10.75 0.51 10.85 ;
      END
   END n_27391

   PIN n_27437
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.35 0.51 48.45 ;
      END
   END n_27437

   PIN n_27439
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.25 0 92.35 0.51 ;
      END
   END n_27439

   PIN n_27513
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.05 295.49 68.15 296 ;
      END
   END n_27513

   PIN n_2774
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 12.45 0 12.55 0.51 ;
      END
   END n_2774

   PIN n_27816
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 107.65 0 107.75 0.51 ;
      END
   END n_27816

   PIN n_27849
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.05 0 20.15 0.51 ;
      END
   END n_27849

   PIN n_27887
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 174.45 0 174.55 0.51 ;
      END
   END n_27887

   PIN n_27899
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 77.45 0 77.55 0.51 ;
      END
   END n_27899

   PIN n_27900
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 152.65 0 152.75 0.51 ;
      END
   END n_27900

   PIN n_27929
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.05 0 104.15 0.51 ;
      END
   END n_27929

   PIN n_27947
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.65 0 41.75 0.51 ;
      END
   END n_27947

   PIN n_27948
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.25 0 104.35 0.51 ;
      END
   END n_27948

   PIN n_28029
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.05 0 102.15 0.51 ;
      END
   END n_28029

   PIN n_28094
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 186.45 0 186.55 0.51 ;
      END
   END n_28094

   PIN n_28111
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.25 0 105.35 0.51 ;
      END
   END n_28111

   PIN n_28189
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.65 0 98.75 0.51 ;
      END
   END n_28189

   PIN n_28201
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 101.45 0 101.55 0.51 ;
      END
   END n_28201

   PIN n_28213
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.05 0 128.15 0.51 ;
      END
   END n_28213

   PIN n_28224
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 191.05 0 191.15 0.51 ;
      END
   END n_28224

   PIN n_28276
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 194.05 0 194.15 0.51 ;
      END
   END n_28276

   PIN n_28296
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 186.25 0 186.35 0.51 ;
      END
   END n_28296

   PIN n_28297
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 190.45 0 190.55 0.51 ;
      END
   END n_28297

   PIN n_28299
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 202.45 0 202.55 0.51 ;
      END
   END n_28299

   PIN n_28326
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 65.05 0 65.15 0.51 ;
      END
   END n_28326

   PIN n_28348
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.45 0 104.55 0.51 ;
      END
   END n_28348

   PIN n_28350
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 114.65 0 114.75 0.51 ;
      END
   END n_28350

   PIN n_28372
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.25 0 185.35 0.51 ;
      END
   END n_28372

   PIN n_28387
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.25 0 116.35 0.51 ;
      END
   END n_28387

   PIN n_28388
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.45 0 116.55 0.51 ;
      END
   END n_28388

   PIN n_28399
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 203.25 0 203.35 0.51 ;
      END
   END n_28399

   PIN n_28430
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.45 0 101.55 0.51 ;
      END
   END n_28430

   PIN n_28431
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 93.45 0 93.55 0.51 ;
      END
   END n_28431

   PIN n_28457
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 184.25 0 184.35 0.51 ;
      END
   END n_28457

   PIN n_28473
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 202.65 0 202.75 0.51 ;
      END
   END n_28473

   PIN n_28474
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.65 0 177.75 0.51 ;
      END
   END n_28474

   PIN n_28500
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 204.05 0 204.15 0.51 ;
      END
   END n_28500

   PIN n_28511
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 93.65 0 93.75 0.51 ;
      END
   END n_28511

   PIN n_28582
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 184.85 0 184.95 0.51 ;
      END
   END n_28582

   PIN n_28583
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 192.85 0 192.95 0.51 ;
      END
   END n_28583

   PIN n_28596
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 207.05 0 207.15 0.51 ;
      END
   END n_28596

   PIN n_28623
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.45 0 103.55 0.51 ;
      END
   END n_28623

   PIN n_28722
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.45 0 92.55 0.51 ;
      END
   END n_28722

   PIN n_28734
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 206.05 0 206.15 0.51 ;
      END
   END n_28734

   PIN n_28743
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 202.25 0 202.35 0.51 ;
      END
   END n_28743

   PIN n_28749
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.45 0 80.55 0.51 ;
      END
   END n_28749

   PIN n_28755
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 194.05 0 194.15 0.51 ;
      END
   END n_28755

   PIN n_28760
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 187.25 0 187.35 0.51 ;
      END
   END n_28760

   PIN n_28763
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 184.45 0 184.55 0.51 ;
      END
   END n_28763

   PIN n_28782
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.65 0 116.75 0.51 ;
      END
   END n_28782

   PIN n_28794
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 21.05 0 21.15 0.51 ;
      END
   END n_28794

   PIN n_28827
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.45 0 128.55 0.51 ;
      END
   END n_28827

   PIN n_28860
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 189.05 0 189.15 0.51 ;
      END
   END n_28860

   PIN n_28864
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.45 0 105.55 0.51 ;
      END
   END n_28864

   PIN n_28869
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.05 0 101.15 0.51 ;
      END
   END n_28869

   PIN n_28888
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.65 0 104.75 0.51 ;
      END
   END n_28888

   PIN n_28929
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 99.25 0 99.35 0.51 ;
      END
   END n_28929

   PIN n_28938
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.65 0 93.75 0.51 ;
      END
   END n_28938

   PIN n_28986
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 115.65 0 115.75 0.51 ;
      END
   END n_28986

   PIN n_29006
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.85 0 100.95 0.51 ;
      END
   END n_29006

   PIN n_29039
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.25 0 115.35 0.51 ;
      END
   END n_29039

   PIN n_29060
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.45 0 114.55 0.51 ;
      END
   END n_29060

   PIN n_29083
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.65 0 102.75 0.51 ;
      END
   END n_29083

   PIN n_29086
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.85 0 96.95 0.51 ;
      END
   END n_29086

   PIN n_29128
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 97.45 0 97.55 0.51 ;
      END
   END n_29128

   PIN n_29133
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 182.65 0 182.75 0.51 ;
      END
   END n_29133

   PIN n_29140
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 183.85 0 183.95 0.51 ;
      END
   END n_29140

   PIN n_29154
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 115.85 0 115.95 0.51 ;
      END
   END n_29154

   PIN n_29251
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.65 0 101.75 0.51 ;
      END
   END n_29251

   PIN n_29269
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.25 0 98.35 0.51 ;
      END
   END n_29269

   PIN n_29329
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 132.45 0 132.55 0.51 ;
      END
   END n_29329

   PIN n_29418
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.85 0 116.95 0.51 ;
      END
   END n_29418

   PIN n_29426
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 117.05 0 117.15 0.51 ;
      END
   END n_29426

   PIN n_29527
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 178.85 0 178.95 0.51 ;
      END
   END n_29527

   PIN n_29608
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.45 0 176.55 0.51 ;
      END
   END n_29608

   PIN n_29625
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 116.05 0 116.15 0.51 ;
      END
   END n_29625

   PIN n_29647
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 170.65 0 170.75 0.51 ;
      END
   END n_29647

   PIN n_29648
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.85 0 92.95 0.51 ;
      END
   END n_29648

   PIN n_29650
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.45 0 93.55 0.51 ;
      END
   END n_29650

   PIN n_29674
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.65 0 91.75 0.51 ;
      END
   END n_29674

   PIN n_29692
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 379.25 0 379.35 0.51 ;
      END
   END n_29692

   PIN n_29701
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.85 0 171.95 0.51 ;
      END
   END n_29701

   PIN n_29719
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.85 0 104.95 0.51 ;
      END
   END n_29719

   PIN n_29721
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.45 0 320.55 0.51 ;
      END
   END n_29721

   PIN n_29723
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 172.65 0 172.75 0.51 ;
      END
   END n_29723

   PIN n_29738
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 175.65 0 175.75 0.51 ;
      END
   END n_29738

   PIN n_29760
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 355.65 0 355.75 0.51 ;
      END
   END n_29760

   PIN n_29815
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 162.85 0 162.95 0.51 ;
      END
   END n_29815

   PIN n_29847
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 99.05 0 99.15 0.51 ;
      END
   END n_29847

   PIN n_29871
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 168.85 0 168.95 0.51 ;
      END
   END n_29871

   PIN n_29888
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 192.25 0 192.35 0.51 ;
      END
   END n_29888

   PIN n_2989
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 51.75 0.51 51.85 ;
      END
   END n_2989

   PIN n_30044
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 334.05 0 334.15 0.51 ;
      END
   END n_30044

   PIN n_3007
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.55 0.51 27.65 ;
      END
   END n_3007

   PIN n_30077
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 370.45 0 370.55 0.51 ;
      END
   END n_30077

   PIN n_30138
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 223.25 0 223.35 0.51 ;
      END
   END n_30138

   PIN n_30169
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 374.05 0 374.15 0.51 ;
      END
   END n_30169

   PIN n_30172
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 335.85 0 335.95 0.51 ;
      END
   END n_30172

   PIN n_30223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 354.85 0 354.95 0.51 ;
      END
   END n_30223

   PIN n_30282
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 372.25 0 372.35 0.51 ;
      END
   END n_30282

   PIN n_30287
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 325.45 0 325.55 0.51 ;
      END
   END n_30287

   PIN n_30333
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.25 0 114.35 0.51 ;
      END
   END n_30333

   PIN n_30356
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 341.85 0 341.95 0.51 ;
      END
   END n_30356

   PIN n_30360
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 403.85 0 403.95 0.51 ;
      END
   END n_30360

   PIN n_30370
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 428.05 0 428.15 0.51 ;
      END
   END n_30370

   PIN n_30373
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 379.85 0 379.95 0.51 ;
      END
   END n_30373

   PIN n_30387
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 375.05 0 375.15 0.51 ;
      END
   END n_30387

   PIN n_30388
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 374.45 0 374.55 0.51 ;
      END
   END n_30388

   PIN n_30391
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 364.85 0 364.95 0.51 ;
      END
   END n_30391

   PIN n_30392
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 363.05 0 363.15 0.51 ;
      END
   END n_30392

   PIN n_30407
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 337.45 0 337.55 0.51 ;
      END
   END n_30407

   PIN n_30426
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 366.25 0 366.35 0.51 ;
      END
   END n_30426

   PIN n_30437
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 391.85 0 391.95 0.51 ;
      END
   END n_30437

   PIN n_30480
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 373.85 0 373.95 0.51 ;
      END
   END n_30480

   PIN n_30487
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 112.45 0 112.55 0.51 ;
      END
   END n_30487

   PIN n_30496
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 127.45 0 127.55 0.51 ;
      END
   END n_30496

   PIN n_30609
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 362.85 0 362.95 0.51 ;
      END
   END n_30609

   PIN n_30616
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 212.65 0 212.75 0.51 ;
      END
   END n_30616

   PIN n_30646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 325.25 0 325.35 0.51 ;
      END
   END n_30646

   PIN n_30656
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 342.25 0 342.35 0.51 ;
      END
   END n_30656

   PIN n_30667
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 361.85 0 361.95 0.51 ;
      END
   END n_30667

   PIN n_30673
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 367.05 0 367.15 0.51 ;
      END
   END n_30673

   PIN n_30685
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 415.85 0 415.95 0.51 ;
      END
   END n_30685

   PIN n_30712
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 333.25 0 333.35 0.51 ;
      END
   END n_30712

   PIN n_30782
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 342.65 0 342.75 0.51 ;
      END
   END n_30782

   PIN n_30795
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 343.25 0 343.35 0.51 ;
      END
   END n_30795

   PIN n_30846
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 364.65 0 364.75 0.51 ;
      END
   END n_30846

   PIN n_30872
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 365.45 0 365.55 0.51 ;
      END
   END n_30872

   PIN n_30945
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 198.85 0 198.95 0.51 ;
      END
   END n_30945

   PIN n_30958
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 356.05 0 356.15 0.51 ;
      END
   END n_30958

   PIN n_30959
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 338.05 0 338.15 0.51 ;
      END
   END n_30959

   PIN n_30977
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 212.25 0 212.35 0.51 ;
      END
   END n_30977

   PIN n_30991
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 331.65 0 331.75 0.51 ;
      END
   END n_30991

   PIN n_31042
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 367.45 0 367.55 0.51 ;
      END
   END n_31042

   PIN n_31076
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 343.45 0 343.55 0.51 ;
      END
   END n_31076

   PIN n_31092
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 346.05 0 346.15 0.51 ;
      END
   END n_31092

   PIN n_31119
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 330.65 0 330.75 0.51 ;
      END
   END n_31119

   PIN n_31120
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 342.4 0 342.6 0.255 ;
      END
   END n_31120

   PIN n_31170
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 344.65 0 344.75 0.51 ;
      END
   END n_31170

   PIN n_31173
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 330.85 0 330.95 0.51 ;
      END
   END n_31173

   PIN n_31184
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 343.05 0 343.15 0.51 ;
      END
   END n_31184

   PIN n_31185
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 342.85 0 342.95 0.51 ;
      END
   END n_31185

   PIN n_31195
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 343.45 0 343.55 0.51 ;
      END
   END n_31195

   PIN n_31218
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 343.65 0 343.75 0.51 ;
      END
   END n_31218

   PIN n_31239
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 360.05 0 360.15 0.51 ;
      END
   END n_31239

   PIN n_31271
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 344.85 0 344.95 0.51 ;
      END
   END n_31271

   PIN n_31355
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 331.05 0 331.15 0.51 ;
      END
   END n_31355

   PIN n_31403
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 340.05 0 340.15 0.51 ;
      END
   END n_31403

   PIN n_31424
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 327.85 0 327.95 0.51 ;
      END
   END n_31424

   PIN n_31460
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 341.65 0 341.75 0.51 ;
      END
   END n_31460

   PIN n_31476
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 361.25 0 361.35 0.51 ;
      END
   END n_31476

   PIN n_31484
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.65 0 126.75 0.51 ;
      END
   END n_31484

   PIN n_31490
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 339.85 0 339.95 0.51 ;
      END
   END n_31490

   PIN n_31494
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 340.05 0 340.15 0.51 ;
      END
   END n_31494

   PIN n_31516
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 357.25 0 357.35 0.51 ;
      END
   END n_31516

   PIN n_3166
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.15 0.51 12.25 ;
      END
   END n_3166

   PIN n_31689
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 351.05 0 351.15 0.51 ;
      END
   END n_31689

   PIN n_31709
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 347.65 0 347.75 0.51 ;
      END
   END n_31709

   PIN n_31727
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 315.85 0 315.95 0.51 ;
      END
   END n_31727

   PIN n_31730
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.05 0 140.15 0.51 ;
      END
   END n_31730

   PIN n_31731
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 59.85 0 59.95 0.51 ;
      END
   END n_31731

   PIN n_31732
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 346.05 0 346.15 0.51 ;
      END
   END n_31732

   PIN n_31734
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 149.05 0 149.15 0.51 ;
      END
   END n_31734

   PIN n_31751
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 307.45 0 307.55 0.51 ;
      END
   END n_31751

   PIN n_31856
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 235.25 0 235.35 0.51 ;
      END
   END n_31856

   PIN n_31919
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 230.45 0 230.55 0.51 ;
      END
   END n_31919

   PIN n_32004
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.45 0 221.55 0.51 ;
      END
   END n_32004

   PIN n_32213
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 216.45 0 216.55 0.51 ;
      END
   END n_32213

   PIN n_32267
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 213.25 0 213.35 0.51 ;
      END
   END n_32267

   PIN n_32307
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 223.85 0 223.95 0.51 ;
      END
   END n_32307

   PIN n_32336
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 214.25 0 214.35 0.51 ;
      END
   END n_32336

   PIN n_32337
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 236.25 0 236.35 0.51 ;
      END
   END n_32337

   PIN n_32344
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.05 0 211.15 0.51 ;
      END
   END n_32344

   PIN n_32386
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.05 0 221.15 0.51 ;
      END
   END n_32386

   PIN n_32387
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 218.65 0 218.75 0.51 ;
      END
   END n_32387

   PIN n_32400
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 130.65 0 130.75 0.51 ;
      END
   END n_32400

   PIN n_32435
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.65 0 224.75 0.51 ;
      END
   END n_32435

   PIN n_32665
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.85 0 163.95 0.51 ;
      END
   END n_32665

   PIN n_32697
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.05 0 164.15 0.51 ;
      END
   END n_32697

   PIN n_32701
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 214.85 0 214.95 0.51 ;
      END
   END n_32701

   PIN n_32779
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.45 0 211.55 0.51 ;
      END
   END n_32779

   PIN n_32785
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.05 0 212.15 0.51 ;
      END
   END n_32785

   PIN n_32805
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 223.25 0 223.35 0.51 ;
      END
   END n_32805

   PIN n_32833
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 236.45 0 236.55 0.51 ;
      END
   END n_32833

   PIN n_32842
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 223.45 0 223.55 0.51 ;
      END
   END n_32842

   PIN n_32845
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 235.85 0 235.95 0.51 ;
      END
   END n_32845

   PIN n_32893
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 222.05 0 222.15 0.51 ;
      END
   END n_32893

   PIN n_32923
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.65 0 151.75 0.51 ;
      END
   END n_32923

   PIN n_32979
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 205.65 0 205.75 0.51 ;
      END
   END n_32979

   PIN n_3304
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.65 0 6.75 0.51 ;
      END
   END n_3304

   PIN n_33066
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 162.85 0 162.95 0.51 ;
      END
   END n_33066

   PIN n_33072
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.25 0 198.35 0.51 ;
      END
   END n_33072

   PIN n_33082
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 235.45 0 235.55 0.51 ;
      END
   END n_33082

   PIN n_33099
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 212.05 0 212.15 0.51 ;
      END
   END n_33099

   PIN n_33111
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.65 0 174.75 0.51 ;
      END
   END n_33111

   PIN n_33201
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 174.65 0 174.75 0.51 ;
      END
   END n_33201

   PIN n_33206
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 186.85 0 186.95 0.51 ;
      END
   END n_33206

   PIN n_33211
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.45 0 198.55 0.51 ;
      END
   END n_33211

   PIN n_33227
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.85 0 198.95 0.51 ;
      END
   END n_33227

   PIN n_33245
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 208.05 0 208.15 0.51 ;
      END
   END n_33245

   PIN n_33253
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 225.45 0 225.55 0.51 ;
      END
   END n_33253

   PIN n_33287
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.45 0 185.55 0.51 ;
      END
   END n_33287

   PIN n_33296
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 213.05 0 213.15 0.51 ;
      END
   END n_33296

   PIN n_33327
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.85 0 220.95 0.51 ;
      END
   END n_33327

   PIN n_33328
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.05 0 199.15 0.51 ;
      END
   END n_33328

   PIN n_33329
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 199.25 0 199.35 0.51 ;
      END
   END n_33329

   PIN n_33422
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.25 0 151.35 0.51 ;
      END
   END n_33422

   PIN n_33463
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 174.85 0 174.95 0.51 ;
      END
   END n_33463

   PIN n_33484
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 252.25 0 252.35 0.51 ;
      END
   END n_33484

   PIN n_3349
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 20.15 0.51 20.25 ;
      END
   END n_3349

   PIN n_33490
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.85 0 151.95 0.51 ;
      END
   END n_33490

   PIN n_33562
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 195.25 0 195.35 0.51 ;
      END
   END n_33562

   PIN n_33566
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 206.45 0 206.55 0.51 ;
      END
   END n_33566

   PIN n_33587
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.65 0 198.75 0.51 ;
      END
   END n_33587

   PIN n_33588
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 201.65 0 201.75 0.51 ;
      END
   END n_33588

   PIN n_33614
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 133.25 0 133.35 0.51 ;
      END
   END n_33614

   PIN n_33630
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.05 0 163.15 0.51 ;
      END
   END n_33630

   PIN n_3365
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 39.55 0.51 39.65 ;
      END
   END n_3365

   PIN n_33653
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 175.05 0 175.15 0.51 ;
      END
   END n_33653

   PIN n_33655
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.85 0 174.95 0.51 ;
      END
   END n_33655

   PIN n_33657
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.25 0 163.35 0.51 ;
      END
   END n_33657

   PIN n_33686
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 452.05 295.49 452.15 296 ;
      END
   END n_33686

   PIN n_33750
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 416.05 0 416.15 0.51 ;
      END
   END n_33750

   PIN n_33757
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 259.85 0 259.95 0.51 ;
      END
   END n_33757

   PIN n_34020
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.65 0 283.75 0.51 ;
      END
   END n_34020

   PIN n_34137
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.25 0 272.35 0.51 ;
      END
   END n_34137

   PIN n_34143
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 286.25 0 286.35 0.51 ;
      END
   END n_34143

   PIN n_34216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.45 0 285.55 0.51 ;
      END
   END n_34216

   PIN n_34299
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.45 0 272.55 0.51 ;
      END
   END n_34299

   PIN n_34438
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 292.05 0 292.15 0.51 ;
      END
   END n_34438

   PIN n_34477
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 283.6 0 283.8 0.255 ;
      END
   END n_34477

   PIN n_34478
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.25 0 199.35 0.51 ;
      END
   END n_34478

   PIN n_34489
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.85 0 284.95 0.51 ;
      END
   END n_34489

   PIN n_34500
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285.05 0 285.15 0.51 ;
      END
   END n_34500

   PIN n_34748
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 298.05 0 298.15 0.51 ;
      END
   END n_34748

   PIN n_34749
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 296.85 0 296.95 0.51 ;
      END
   END n_34749

   PIN n_34758
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.05 0 281.15 0.51 ;
      END
   END n_34758

   PIN n_34759
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 283.25 0 283.35 0.51 ;
      END
   END n_34759

   PIN n_34760
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 288.25 0 288.35 0.51 ;
      END
   END n_34760

   PIN n_34775
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 286.45 0 286.55 0.51 ;
      END
   END n_34775

   PIN n_34788
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.65 0 271.75 0.51 ;
      END
   END n_34788

   PIN n_3487
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 18.95 0.51 19.05 ;
      END
   END n_3487

   PIN n_34902
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 287.65 0 287.75 0.51 ;
      END
   END n_34902

   PIN n_34904
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 295.45 0 295.55 0.51 ;
      END
   END n_34904

   PIN n_34943
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.65 0 291.75 0.51 ;
      END
   END n_34943

   PIN n_35025
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.85 0 294.95 0.51 ;
      END
   END n_35025

   PIN n_35036
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.85 0 292.95 0.51 ;
      END
   END n_35036

   PIN n_35105
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.65 0 294.75 0.51 ;
      END
   END n_35105

   PIN n_35129
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.25 0 285.35 0.51 ;
      END
   END n_35129

   PIN n_35131
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 280.45 0 280.55 0.51 ;
      END
   END n_35131

   PIN n_35134
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.45 0 292.55 0.51 ;
      END
   END n_35134

   PIN n_35140
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.25 0 283.35 0.51 ;
      END
   END n_35140

   PIN n_35143
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 286.65 0 286.75 0.51 ;
      END
   END n_35143

   PIN n_35375
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 272.25 0 272.35 0.51 ;
      END
   END n_35375

   PIN n_35580
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 296.25 0 296.35 0.51 ;
      END
   END n_35580

   PIN n_4090
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.55 0.51 32.65 ;
      END
   END n_4090

   PIN n_4133
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.65 0 20.75 0.51 ;
      END
   END n_4133

   PIN n_4333
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.25 0 4.35 0.51 ;
      END
   END n_4333

   PIN n_4413
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.25 0 33.35 0.51 ;
      END
   END n_4413

   PIN n_4526
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 19.15 0.51 19.25 ;
      END
   END n_4526

   PIN n_4634
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 244.55 0.51 244.65 ;
      END
   END n_4634

   PIN n_4673
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 100.35 0.51 100.45 ;
      END
   END n_4673

   PIN n_4761
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.35 0.51 12.45 ;
      END
   END n_4761

   PIN n_4889
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 19.35 0.51 19.45 ;
      END
   END n_4889

   PIN n_4902
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 267.95 0.51 268.05 ;
      END
   END n_4902

   PIN n_4922
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.35 0.51 64.45 ;
      END
   END n_4922

   PIN n_5077
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 20.35 0.51 20.45 ;
      END
   END n_5077

   PIN n_62095
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.35 0.51 26.45 ;
      END
   END n_62095

   PIN n_63235
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.95 0.51 30.05 ;
      END
   END n_63235

   PIN n_63270
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.75 0.51 32.85 ;
      END
   END n_63270

   PIN n_63281
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.85 0 21.95 0.51 ;
      END
   END n_63281

   PIN n_63816
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.45 0 77.55 0.51 ;
      END
   END n_63816

   PIN n_64050
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.05 0 74.15 0.51 ;
      END
   END n_64050

   PIN n_64089
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 76.25 0 76.35 0.51 ;
      END
   END n_64089

   PIN n_64141
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 75.45 0 75.55 0.51 ;
      END
   END n_64141

   PIN n_64164
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.65 0 80.75 0.51 ;
      END
   END n_64164

   PIN n_64228
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.85 0 72.95 0.51 ;
      END
   END n_64228

   PIN n_64301
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 66.05 0 66.15 0.51 ;
      END
   END n_64301

   PIN n_64325
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 63.85 0 63.95 0.51 ;
      END
   END n_64325

   PIN n_64384
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 74.85 0 74.95 0.51 ;
      END
   END n_64384

   PIN n_64437
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.25 0 74.35 0.51 ;
      END
   END n_64437

   PIN n_64570
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.85 0 68.95 0.51 ;
      END
   END n_64570

   PIN n_64704
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.85 0 80.95 0.51 ;
      END
   END n_64704

   PIN n_64735
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 73.45 0 73.55 0.51 ;
      END
   END n_64735

   PIN n_64770
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 136.35 0.51 136.45 ;
      END
   END n_64770

   PIN n_64800
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.65 0 67.75 0.51 ;
      END
   END n_64800

   PIN n_64801
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 63.25 0 63.35 0.51 ;
      END
   END n_64801

   PIN n_64811
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 196.75 0.51 196.85 ;
      END
   END n_64811

   PIN n_64946
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 62.05 0 62.15 0.51 ;
      END
   END n_64946

   PIN n_64982
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 60.25 0 60.35 0.51 ;
      END
   END n_64982

   PIN n_65063
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 60.45 0 60.55 0.51 ;
      END
   END n_65063

   PIN n_65156
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.45 0 64.55 0.51 ;
      END
   END n_65156

   PIN n_65198
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 63.65 0 63.75 0.51 ;
      END
   END n_65198

   PIN n_65585
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.05 0 85.15 0.51 ;
      END
   END n_65585

   PIN n_65644
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 11.75 0.51 11.85 ;
      END
   END n_65644

   PIN n_65659
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.85 295.49 163.95 296 ;
      END
   END n_65659

   PIN n_65667
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.25 0 81.35 0.51 ;
      END
   END n_65667

   PIN n_65746
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 11.95 0.51 12.05 ;
      END
   END n_65746

   PIN n_65780
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 47.05 0 47.15 0.51 ;
      END
   END n_65780

   PIN n_65811
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 10.15 0.51 10.25 ;
      END
   END n_65811

   PIN n_65824
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 52.05 0 52.15 0.51 ;
      END
   END n_65824

   PIN n_65827
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.05 295.49 164.15 296 ;
      END
   END n_65827

   PIN n_65830
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.55 0.51 39.65 ;
      END
   END n_65830

   PIN n_65889
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.35 0.51 123.45 ;
      END
   END n_65889

   PIN n_65900
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 87.25 0 87.35 0.51 ;
      END
   END n_65900

   PIN n_65921
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 83.65 0 83.75 0.51 ;
      END
   END n_65921

   PIN n_65938
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 47.45 0 47.55 0.51 ;
      END
   END n_65938

   PIN n_65939
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44.85 0 44.95 0.51 ;
      END
   END n_65939

   PIN n_65940
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.55 0.51 32.65 ;
      END
   END n_65940

   PIN n_65963
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 87.65 0 87.75 0.51 ;
      END
   END n_65963

   PIN n_66043
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 46.25 0 46.35 0.51 ;
      END
   END n_66043

   PIN n_66049
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44.65 0 44.75 0.51 ;
      END
   END n_66049

   PIN n_66062
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.95 0.51 39.05 ;
      END
   END n_66062

   PIN n_66063
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.75 0.51 112.85 ;
      END
   END n_66063

   PIN n_66064
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.55 0.51 111.65 ;
      END
   END n_66064

   PIN n_66072
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 86.65 0 86.75 0.51 ;
      END
   END n_66072

   PIN n_66147
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.85 0 36.95 0.51 ;
      END
   END n_66147

   PIN n_66148
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 46.45 0 46.55 0.51 ;
      END
   END n_66148

   PIN n_66150
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 82.65 0 82.75 0.51 ;
      END
   END n_66150

   PIN n_66151
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.65 0 92.75 0.51 ;
      END
   END n_66151

   PIN n_66163
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.95 0.51 29.05 ;
      END
   END n_66163

   PIN n_66220
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 79.25 0 79.35 0.51 ;
      END
   END n_66220

   PIN n_66234
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.15 0.51 32.25 ;
      END
   END n_66234

   PIN n_66256
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 86.05 0 86.15 0.51 ;
      END
   END n_66256

   PIN n_66277
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.75 0.51 39.85 ;
      END
   END n_66277

   PIN n_66320
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.05 295.49 80.15 296 ;
      END
   END n_66320

   PIN n_66322
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 84.85 0 84.95 0.51 ;
      END
   END n_66322

   PIN n_66366
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.35 0.51 111.45 ;
      END
   END n_66366

   PIN n_66379
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 12.15 0.51 12.25 ;
      END
   END n_66379

   PIN n_66409
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.25 0 88.35 0.51 ;
      END
   END n_66409

   PIN n_66421
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.95 0.51 40.05 ;
      END
   END n_66421

   PIN n_66434
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.15 0.51 40.25 ;
      END
   END n_66434

   PIN n_66456
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.65 0 78.75 0.51 ;
      END
   END n_66456

   PIN n_66462
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 23.15 0.51 23.25 ;
      END
   END n_66462

   PIN n_66488
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.75 0.51 37.85 ;
      END
   END n_66488

   PIN n_66520
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 22.8 0 23 0.255 ;
      END
   END n_66520

   PIN n_66544
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.85 0 40.95 0.51 ;
      END
   END n_66544

   PIN n_66548
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.05 0 80.15 0.51 ;
      END
   END n_66548

   PIN n_66565
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 21.85 0 21.95 0.51 ;
      END
   END n_66565

   PIN n_66570
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 27.75 0.51 27.85 ;
      END
   END n_66570

   PIN n_66577
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.35 0.51 38.45 ;
      END
   END n_66577

   PIN n_66582
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 87.65 0 87.75 0.51 ;
      END
   END n_66582

   PIN n_66586
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 22.05 0 22.15 0.51 ;
      END
   END n_66586

   PIN n_66593
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 81.85 0 81.95 0.51 ;
      END
   END n_66593

   PIN n_66595
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44.25 0 44.35 0.51 ;
      END
   END n_66595

   PIN n_66622
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.35 0.51 40.45 ;
      END
   END n_66622

   PIN n_66638
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 22.25 0 22.35 0.51 ;
      END
   END n_66638

   PIN n_66647
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 45.25 0 45.35 0.51 ;
      END
   END n_66647

   PIN n_66650
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.85 0 83.95 0.51 ;
      END
   END n_66650

   PIN n_66655
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.95 0.51 113.05 ;
      END
   END n_66655

   PIN n_66706
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 19.55 0.51 19.65 ;
      END
   END n_66706

   PIN n_66765
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 39.75 0.51 39.85 ;
      END
   END n_66765

   PIN n_66766
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.55 0.51 34.65 ;
      END
   END n_66766

   PIN n_66777
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 85.05 0 85.15 0.51 ;
      END
   END n_66777

   PIN n_66845
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 38.65 0 38.75 0.51 ;
      END
   END n_66845

   PIN n_66858
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.25 0 80.35 0.51 ;
      END
   END n_66858

   PIN n_66866
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 135.95 0.51 136.05 ;
      END
   END n_66866

   PIN n_66877
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.95 0.51 38.05 ;
      END
   END n_66877

   PIN n_66939
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 136.15 0.51 136.25 ;
      END
   END n_66939

   PIN n_66996
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 66.25 0 66.35 0.51 ;
      END
   END n_66996

   PIN n_67014
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 82.05 0 82.15 0.51 ;
      END
   END n_67014

   PIN n_67059
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 41.05 0 41.15 0.51 ;
      END
   END n_67059

   PIN n_67072
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.25 0 36.35 0.51 ;
      END
   END n_67072

   PIN n_67086
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 39.95 0.51 40.05 ;
      END
   END n_67086

   PIN n_67110
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.55 0.51 123.65 ;
      END
   END n_67110

   PIN n_67204
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 13.25 0 13.35 0.51 ;
      END
   END n_67204

   PIN n_67239
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.65 0 10.75 0.51 ;
      END
   END n_67239

   PIN n_67252
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 0.65 0 0.75 0.51 ;
      END
   END n_67252

   PIN n_67253
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 35.45 0 35.55 0.51 ;
      END
   END n_67253

   PIN n_67287
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.55 0.51 64.65 ;
      END
   END n_67287

   PIN n_6732
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 167.45 0 167.55 0.51 ;
      END
   END n_6732

   PIN n_67320
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 42.65 0 42.75 0.51 ;
      END
   END n_67320

   PIN n_67524
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 46.05 0 46.15 0.51 ;
      END
   END n_67524

   PIN n_67561
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.05 0 57.15 0.51 ;
      END
   END n_67561

   PIN n_67606
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 92.85 0 92.95 0.51 ;
      END
   END n_67606

   PIN n_67801
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.45 0 55.55 0.51 ;
      END
   END n_67801

   PIN n_67898
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 81.05 0 81.15 0.51 ;
      END
   END n_67898

   PIN n_67995
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.45 0 57.55 0.51 ;
      END
   END n_67995

   PIN n_68021
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 54.05 0 54.15 0.51 ;
      END
   END n_68021

   PIN n_68043
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 53.05 0 53.15 0.51 ;
      END
   END n_68043

   PIN n_68092
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.85 0 50.95 0.51 ;
      END
   END n_68092

   PIN n_68186
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.65 0 55.75 0.51 ;
      END
   END n_68186

   PIN n_68213
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 65.85 0 65.95 0.51 ;
      END
   END n_68213

   PIN n_68361
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.45 0 56.55 0.51 ;
      END
   END n_68361

   PIN n_68364
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.65 0 59.75 0.51 ;
      END
   END n_68364

   PIN n_68492
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 54.45 0 54.55 0.51 ;
      END
   END n_68492

   PIN n_68493
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 53.85 0 53.95 0.51 ;
      END
   END n_68493

   PIN n_68509
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 53.65 0 53.75 0.51 ;
      END
   END n_68509

   PIN n_68549
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.65 0 57.75 0.51 ;
      END
   END n_68549

   PIN n_68730
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 93.85 0 93.95 0.51 ;
      END
   END n_68730

   PIN n_68839
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 53.25 0 53.35 0.51 ;
      END
   END n_68839

   PIN n_68842
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 53.45 0 53.55 0.51 ;
      END
   END n_68842

   PIN n_69233
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 39.45 0 39.55 0.51 ;
      END
   END n_69233

   PIN n_69250
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.25 0 24.35 0.51 ;
      END
   END n_69250

   PIN n_69476
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 342.05 0 342.15 0.51 ;
      END
   END n_69476

   PIN n_69494
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 64.85 0 64.95 0.51 ;
      END
   END n_69494

   PIN n_69523
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.45 0 307.55 0.51 ;
      END
   END n_69523

   PIN n_69725
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 332.85 0 332.95 0.51 ;
      END
   END n_69725

   PIN n_69742
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 73.05 0 73.15 0.51 ;
      END
   END n_69742

   PIN n_69765
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 331.45 0 331.55 0.51 ;
      END
   END n_69765

   PIN n_69846
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.05 0 307.15 0.51 ;
      END
   END n_69846

   PIN n_69856
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.65 0 72.75 0.51 ;
      END
   END n_69856

   PIN n_69945
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37.25 0 37.35 0.51 ;
      END
   END n_69945

   PIN n_70024
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.85 0 63.95 0.51 ;
      END
   END n_70024

   PIN n_70049
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.45 0 36.55 0.51 ;
      END
   END n_70049

   PIN n_70182
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.45 0 318.55 0.51 ;
      END
   END n_70182

   PIN n_70208
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37.45 0 37.55 0.51 ;
      END
   END n_70208

   PIN n_70223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 307.65 0 307.75 0.51 ;
      END
   END n_70223

   PIN n_70238
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 43.65 0 43.75 0.51 ;
      END
   END n_70238

   PIN n_70269
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.65 0 320.75 0.51 ;
      END
   END n_70269

   PIN n_70323
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.65 0 320.75 0.51 ;
      END
   END n_70323

   PIN n_70327
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.85 0 318.95 0.51 ;
      END
   END n_70327

   PIN n_70356
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 295.05 0 295.15 0.51 ;
      END
   END n_70356

   PIN n_70391
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.25 0 307.35 0.51 ;
      END
   END n_70391

   PIN n_70403
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 332.4 0 332.6 0.255 ;
      END
   END n_70403

   PIN n_70473
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.05 0 319.15 0.51 ;
      END
   END n_70473

   PIN n_70483
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.85 0 320.95 0.51 ;
      END
   END n_70483

   PIN n_70489
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.05 0 319.15 0.51 ;
      END
   END n_70489

   PIN n_70532
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.25 0 319.35 0.51 ;
      END
   END n_70532

   PIN n_70542
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.85 0 320.95 0.51 ;
      END
   END n_70542

   PIN n_70558
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 65.45 0 65.55 0.51 ;
      END
   END n_70558

   PIN n_70643
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 313.05 0 313.15 0.51 ;
      END
   END n_70643

   PIN n_70646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 43.85 0 43.95 0.51 ;
      END
   END n_70646

   PIN n_70748
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 307.85 0 307.95 0.51 ;
      END
   END n_70748

   PIN n_70793
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.85 0 306.95 0.51 ;
      END
   END n_70793

   PIN n_70794
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.05 0 308.15 0.51 ;
      END
   END n_70794

   PIN n_70803
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 67.45 0 67.55 0.51 ;
      END
   END n_70803

   PIN n_70857
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 296.45 0 296.55 0.51 ;
      END
   END n_70857

   PIN n_70928
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.25 0 308.35 0.51 ;
      END
   END n_70928

   PIN n_70933
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.05 0 321.15 0.51 ;
      END
   END n_70933

   PIN n_71006
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.25 0 321.35 0.51 ;
      END
   END n_71006

   PIN n_71030
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.45 0 308.55 0.51 ;
      END
   END n_71030

   PIN n_71082
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.65 0 307.75 0.51 ;
      END
   END n_71082

   PIN n_71149
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.95 0.51 69.05 ;
      END
   END n_71149

   PIN n_71253
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.95 0.51 59.05 ;
      END
   END n_71253

   PIN n_71285
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.85 0 56.95 0.51 ;
      END
   END n_71285

   PIN n_71297
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.45 0 78.55 0.51 ;
      END
   END n_71297

   PIN n_738
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.45 0 18.55 0.51 ;
      END
   END n_738

   PIN n_75924
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 51.95 0.51 52.05 ;
      END
   END n_75924

   PIN n_75925
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.65 0 28.75 0.51 ;
      END
   END n_75925

   PIN n_76109
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.25 0 56.35 0.51 ;
      END
   END n_76109

   PIN n_76206
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 36.35 0.51 36.45 ;
      END
   END n_76206

   PIN n_76260
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 76.2 0 76.4 0.255 ;
      END
   END n_76260

   PIN n_76261
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 26.25 0 26.35 0.51 ;
      END
   END n_76261

   PIN n_76271
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 23.35 0.51 23.45 ;
      END
   END n_76271

   PIN n_76280
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.45 0 56.55 0.51 ;
      END
   END n_76280

   PIN n_76281
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 49.95 0.51 50.05 ;
      END
   END n_76281

   PIN n_76282
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 40.15 0.51 40.25 ;
      END
   END n_76282

   PIN n_76283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 27.25 0 27.35 0.51 ;
      END
   END n_76283

   PIN n_76292
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 40.25 0 40.35 0.51 ;
      END
   END n_76292

   PIN n_76347
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.45 0 29.55 0.51 ;
      END
   END n_76347

   PIN n_76417
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.85 0 33.95 0.51 ;
      END
   END n_76417

   PIN n_76638
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 27.05 0 27.15 0.51 ;
      END
   END n_76638

   PIN n_76852
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 25.05 0 25.15 0.51 ;
      END
   END n_76852

   PIN n_76965
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 52.15 0.51 52.25 ;
      END
   END n_76965

   PIN n_77013
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 30.65 0 30.75 0.51 ;
      END
   END n_77013

   PIN n_77047
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.45 0 25.55 0.51 ;
      END
   END n_77047

   PIN n_77053
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 63.55 0.51 63.65 ;
      END
   END n_77053

   PIN n_77442
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.05 0 25.15 0.51 ;
      END
   END n_77442

   PIN n_77600
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.15 0.51 77.25 ;
      END
   END n_77600

   PIN n_78116
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.65 0 31.75 0.51 ;
      END
   END n_78116

   PIN n_823
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.95 0.51 42.05 ;
      END
   END n_823

   PIN n_923
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.25 0 25.35 0.51 ;
      END
   END n_923

   PIN u0_L7_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.25 0 128.35 0.51 ;
      END
   END u0_L7_13_

   PIN u0_L7_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.25 0 140.35 0.51 ;
      END
   END u0_L7_3_

   PIN u0_L7_reg_14__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 118.05 0 118.15 0.51 ;
      END
   END u0_L7_reg_14__Q

   PIN u0_L7_reg_17__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 116.25 0 116.35 0.51 ;
      END
   END u0_L7_reg_17__Q

   PIN u0_L7_reg_18__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 275.45 0 275.55 0.51 ;
      END
   END u0_L7_reg_18__Q

   PIN u0_L8_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.45 0 197.55 0.51 ;
      END
   END u0_L8_12_

   PIN u0_L8_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.65 0 119.75 0.51 ;
      END
   END u0_L8_28_

   PIN u0_L8_reg_7__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 235.85 0 235.95 0.51 ;
      END
   END u0_L8_reg_7__Q

   PIN u0_L9_26_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 192.65 0 192.75 0.51 ;
      END
   END u0_L9_26_

   PIN u0_R10_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 548.69 11.15 549.2 11.25 ;
      END
   END u0_R10_23_

   PIN u0_R3_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 37.55 0.51 37.65 ;
      END
   END u0_R3_11_

   PIN u0_R4_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 62.55 0.51 62.65 ;
      END
   END u0_R4_1_

   PIN u0_R5_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 1.45 0 1.55 0.51 ;
      END
   END u0_R5_11_

   PIN u0_R5_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 25.65 0 25.75 0.51 ;
      END
   END u0_R5_14_

   PIN u0_R5_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.65 0 38.75 0.51 ;
      END
   END u0_R5_15_

   PIN u0_R5_19_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 18.65 0 18.75 0.51 ;
      END
   END u0_R5_19_

   PIN u0_R5_29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.65 0 138.75 0.51 ;
      END
   END u0_R5_29_

   PIN u0_R6_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 129.25 0 129.35 0.51 ;
      END
   END u0_R6_13_

   PIN u0_R6_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 40.85 0 40.95 0.51 ;
      END
   END u0_R6_1_

   PIN u0_R6_20_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 105.05 0 105.15 0.51 ;
      END
   END u0_R6_20_

   PIN u0_R6_30_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 94.05 0 94.15 0.51 ;
      END
   END u0_R6_30_

   PIN u0_R6_31_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 52.45 0 52.55 0.51 ;
      END
   END u0_R6_31_

   PIN u0_R6_32_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 52.65 0 52.75 0.51 ;
      END
   END u0_R6_32_

   PIN u0_R7_17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 58.45 0 58.55 0.51 ;
      END
   END u0_R7_17_

   PIN u0_R7_19_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 190.85 0 190.95 0.51 ;
      END
   END u0_R7_19_

   PIN u0_R7_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 112.25 0 112.35 0.51 ;
      END
   END u0_R7_7_

   PIN u0_R8_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.25 0 138.35 0.51 ;
      END
   END u0_R8_12_

   PIN u0_R8_17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.65 0 308.75 0.51 ;
      END
   END u0_R8_17_

   PIN u0_R8_20_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 83.45 0 83.55 0.51 ;
      END
   END u0_R8_20_

   PIN u0_R8_26_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 295.45 0 295.55 0.51 ;
      END
   END u0_R8_26_

   PIN u0_R8_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.05 0 260.15 0.51 ;
      END
   END u0_R8_3_

   PIN u0_R8_9_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 311.05 0 311.15 0.51 ;
      END
   END u0_R8_9_

   PIN u0_R9_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 440.05 0 440.15 0.51 ;
      END
   END u0_R9_12_

   PIN u0_R9_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 204.85 0 204.95 0.51 ;
      END
   END u0_R9_1_

   PIN u0_key_r_55_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 42.85 0 42.95 0.51 ;
      END
   END u0_key_r_55_

   PIN u0_uk_K_r_239
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 78.25 0 78.35 0.51 ;
      END
   END u0_uk_K_r_239

   PIN u0_uk_K_r_264
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 20.35 0.51 20.45 ;
      END
   END u0_uk_K_r_264

   PIN u0_uk_K_r_349
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 43.05 0 43.15 0.51 ;
      END
   END u0_uk_K_r_349

   PIN u0_uk_K_r_353
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 9.25 0 9.35 0.51 ;
      END
   END u0_uk_K_r_353

   PIN u0_uk_K_r_361
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.65 0 16.75 0.51 ;
      END
   END u0_uk_K_r_361

   PIN u0_uk_K_r_373
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 20.95 0.51 21.05 ;
      END
   END u0_uk_K_r_373

   PIN u0_uk_K_r_383
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 24.05 0 24.15 0.51 ;
      END
   END u0_uk_K_r_383

   PIN u0_uk_K_r_387
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.75 0.51 34.85 ;
      END
   END u0_uk_K_r_387

   PIN u0_uk_K_r_390
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.75 0.51 27.85 ;
      END
   END u0_uk_K_r_390

   PIN u0_uk_K_r_399
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.75 0.51 26.85 ;
      END
   END u0_uk_K_r_399

   PIN u0_uk_K_r_412
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.65 0 36.75 0.51 ;
      END
   END u0_uk_K_r_412

   PIN u0_uk_K_r_433
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.85 0 12.95 0.51 ;
      END
   END u0_uk_K_r_433

   PIN u0_uk_K_r_436
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.05 0 16.15 0.51 ;
      END
   END u0_uk_K_r_436

   PIN u0_uk_K_r_463
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 37.75 0.51 37.85 ;
      END
   END u0_uk_K_r_463

   PIN u0_uk_K_r_469
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.85 0 10.95 0.51 ;
      END
   END u0_uk_K_r_469

   PIN u0_uk_K_r_492
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.05 0 12.15 0.51 ;
      END
   END u0_uk_K_r_492

   PIN u0_uk_K_r_518
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 25.45 0 25.55 0.51 ;
      END
   END u0_uk_K_r_518

   PIN u0_uk_K_r_523
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 52.35 0.51 52.45 ;
      END
   END u0_uk_K_r_523

   PIN u0_uk_K_r_547
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 14.65 0 14.75 0.51 ;
      END
   END u0_uk_K_r_547

   PIN u1_IP_22_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 76.45 0 76.55 0.51 ;
      END
   END u1_IP_22_

   PIN u1_L11_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.25 0 319.35 0.51 ;
      END
   END u1_L11_7_

   PIN u1_R10_29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.95 0.51 41.05 ;
      END
   END u1_R10_29_

   PIN u1_R10_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 24.55 0.51 24.65 ;
      END
   END u1_R10_4_

   PIN u1_desIn_r_reg_28__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 92.05 0 92.15 0.51 ;
      END
   END u1_desIn_r_reg_28__Q

   PIN u1_desIn_r_reg_54__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 58.05 0 58.15 0.51 ;
      END
   END u1_desIn_r_reg_54__Q

   PIN u2_L7_reg_12__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 392.05 0 392.15 0.51 ;
      END
   END u2_L7_reg_12__Q

   PIN u2_L7_reg_7__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 366.85 0 366.95 0.51 ;
      END
   END u2_L7_reg_7__Q

   PIN FE_OFN1018_n_6197
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 37.65 0 37.75 0.51 ;
      END
   END FE_OFN1018_n_6197

   PIN FE_OFN1021_n_3701
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 3.45 0 3.55 0.51 ;
      END
   END FE_OFN1021_n_3701

   PIN FE_OFN1068_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.05 0 28.15 0.51 ;
      END
   END FE_OFN1068_n_116

   PIN FE_OFN1094_g303299_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 4.65 0 4.75 0.51 ;
      END
   END FE_OFN1094_g303299_p

   PIN FE_OFN1105_n_6021
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.25 0 59.35 0.51 ;
      END
   END FE_OFN1105_n_6021

   PIN FE_OFN1224_n_6583
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 83.85 0 83.95 0.51 ;
      END
   END FE_OFN1224_n_6583

   PIN FE_OFN1292_n_4098
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.85 0 23.95 0.51 ;
      END
   END FE_OFN1292_n_4098

   PIN FE_OFN1338_n_117596
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.45 0 199.55 0.51 ;
      END
   END FE_OFN1338_n_117596

   PIN FE_OFN1381_n_6875
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.65 0 159.75 0.51 ;
      END
   END FE_OFN1381_n_6875

   PIN FE_OFN1578_n_3047
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.85 0 6.95 0.51 ;
      END
   END FE_OFN1578_n_3047

   PIN FE_OFN1646_n_6731
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 169.05 0 169.15 0.51 ;
      END
   END FE_OFN1646_n_6731

   PIN FE_OFN1735_n_64033
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 88.7 0.255 88.9 ;
      END
   END FE_OFN1735_n_64033

   PIN FE_OFN1933_n_69492
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 77.85 0 77.95 0.51 ;
      END
   END FE_OFN1933_n_69492

   PIN FE_OFN1958_n_6873
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 94.65 0 94.75 0.51 ;
      END
   END FE_OFN1958_n_6873

   PIN FE_OFN2009_n_27918
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 57.65 0 57.75 0.51 ;
      END
   END FE_OFN2009_n_27918

   PIN FE_OFN2013_n_23906
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.45 0 12.55 0.51 ;
      END
   END FE_OFN2013_n_23906

   PIN FE_OFN2114_n_19614
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.65 0 56.75 0.51 ;
      END
   END FE_OFN2114_n_19614

   PIN FE_OFN2221_g302057_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.05 0 3.15 0.51 ;
      END
   END FE_OFN2221_g302057_p

   PIN FE_OFN2276_n_27867
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.85 0 34.95 0.51 ;
      END
   END FE_OFN2276_n_27867

   PIN FE_OFN2316_n_65154
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.85 0 64.95 0.51 ;
      END
   END FE_OFN2316_n_65154

   PIN FE_OFN2333_n_23919
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 11.35 0.51 11.45 ;
      END
   END FE_OFN2333_n_23919

   PIN FE_OFN2351_n_27890
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.45 0 27.55 0.51 ;
      END
   END FE_OFN2351_n_27890

   PIN FE_OFN2406_n_13312
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 1.65 0 1.75 0.51 ;
      END
   END FE_OFN2406_n_13312

   PIN FE_OFN2417_n_26365
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 172.15 0.51 172.25 ;
      END
   END FE_OFN2417_n_26365

   PIN FE_OFN2472_n_117820
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 18.45 0 18.55 0.51 ;
      END
   END FE_OFN2472_n_117820

   PIN FE_OFN2503_n_5437
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.25 0 77.35 0.51 ;
      END
   END FE_OFN2503_n_5437

   PIN FE_OFN2504_n_4918
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.05 0 8.15 0.51 ;
      END
   END FE_OFN2504_n_4918

   PIN FE_OFN2537_n_65517
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.85 0 7.95 0.51 ;
      END
   END FE_OFN2537_n_65517

   PIN FE_OFN2677_n_23958
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.45 0 42.55 0.51 ;
      END
   END FE_OFN2677_n_23958

   PIN FE_OFN2719_n_25980
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 25.25 0 25.35 0.51 ;
      END
   END FE_OFN2719_n_25980

   PIN FE_OFN2786_n_5684
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.85 0 36.95 0.51 ;
      END
   END FE_OFN2786_n_5684

   PIN FE_OFN2930_n_4064
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15.85 0 15.95 0.51 ;
      END
   END FE_OFN2930_n_4064

   PIN FE_OFN2965_n_4653
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.05 0 19.15 0.51 ;
      END
   END FE_OFN2965_n_4653

   PIN FE_OFN2975_n_65768
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 3.25 0 3.35 0.51 ;
      END
   END FE_OFN2975_n_65768

   PIN FE_OFN2982_n_65436
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.85 0 43.95 0.51 ;
      END
   END FE_OFN2982_n_65436

   PIN FE_OFN2993_n_6198
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15.25 0 15.35 0.51 ;
      END
   END FE_OFN2993_n_6198

   PIN FE_OFN3017_n_69766
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 78.85 0 78.95 0.51 ;
      END
   END FE_OFN3017_n_69766

   PIN FE_OFN3049_n_3016
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.25 0 27.35 0.51 ;
      END
   END FE_OFN3049_n_3016

   PIN FE_OFN3146_n_35477
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.85 0 282.95 0.51 ;
      END
   END FE_OFN3146_n_35477

   PIN FE_OFN3152_n_25832
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.45 0 36.55 0.51 ;
      END
   END FE_OFN3152_n_25832

   PIN FE_OFN3164_n_2780
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.05 0 24.15 0.51 ;
      END
   END FE_OFN3164_n_2780

   PIN FE_OFN3226_g302039_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.05 0 14.15 0.51 ;
      END
   END FE_OFN3226_g302039_p

   PIN FE_OFN3240_n_4790
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.55 0.51 26.65 ;
      END
   END FE_OFN3240_n_4790

   PIN FE_OFN324_n_70684
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 332.45 0 332.55 0.51 ;
      END
   END FE_OFN324_n_70684

   PIN FE_OFN326_n_70685
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.05 0 320.15 0.51 ;
      END
   END FE_OFN326_n_70685

   PIN FE_OFN3278_n_39
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.85 0 3.95 0.51 ;
      END
   END FE_OFN3278_n_39

   PIN FE_OFN3318_n_500
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 99 295.745 99.2 296 ;
      END
   END FE_OFN3318_n_500

   PIN FE_OFN3319_n_500
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.9 0.255 96.1 ;
      END
   END FE_OFN3319_n_500

   PIN FE_OFN3365_n_5443
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.05 0 20.15 0.51 ;
      END
   END FE_OFN3365_n_5443

   PIN FE_OFN3399_n_7096
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.85 0 6.95 0.51 ;
      END
   END FE_OFN3399_n_7096

   PIN FE_OFN3463_n_67106
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.75 0.51 41.85 ;
      END
   END FE_OFN3463_n_67106

   PIN FE_OFN3485_n_1596
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.45 0 11.55 0.51 ;
      END
   END FE_OFN3485_n_1596

   PIN FE_OFN3516_n_23820
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 19.75 0.51 19.85 ;
      END
   END FE_OFN3516_n_23820

   PIN FE_OFN3542_g302047_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.85 0 5.95 0.51 ;
      END
   END FE_OFN3542_g302047_p

   PIN FE_OFN3627_n_4557
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.65 0 33.75 0.51 ;
      END
   END FE_OFN3627_n_4557

   PIN FE_OFN373_n_66358
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 37.25 0 37.35 0.51 ;
      END
   END FE_OFN373_n_66358

   PIN FE_OFN375_n_65823
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 22.45 0 22.55 0.51 ;
      END
   END FE_OFN375_n_65823

   PIN FE_OFN3784_n_60
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.15 0.51 27.25 ;
      END
   END FE_OFN3784_n_60

   PIN FE_OFN3799_n_23840
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.35 0.51 16.45 ;
      END
   END FE_OFN3799_n_23840

   PIN FE_OFN3858_n_68782
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 53.25 0 53.35 0.51 ;
      END
   END FE_OFN3858_n_68782

   PIN FE_OFN3909_n_5532
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 14.85 0 14.95 0.51 ;
      END
   END FE_OFN3909_n_5532

   PIN FE_OFN3914_n_29934
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 362.45 0 362.55 0.51 ;
      END
   END FE_OFN3914_n_29934

   PIN FE_OFN3965_n_9884
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.15 0.51 34.25 ;
      END
   END FE_OFN3965_n_9884

   PIN FE_OFN4124_g302043_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 4.85 0 4.95 0.51 ;
      END
   END FE_OFN4124_g302043_p

   PIN FE_OFN4143_n_29936
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.45 0 140.55 0.51 ;
      END
   END FE_OFN4143_n_29936

   PIN FE_OFN4244_n_29500
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 178.05 0 178.15 0.51 ;
      END
   END FE_OFN4244_n_29500

   PIN FE_OFN4315_n_104
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 32.6 0 32.8 0.255 ;
      END
   END FE_OFN4315_n_104

   PIN FE_OFN4359_n_20
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 23.2 0 23.4 0.255 ;
      END
   END FE_OFN4359_n_20

   PIN FE_OFN4412_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.3 0.255 24.5 ;
      END
   END FE_OFN4412_decrypt

   PIN FE_OFN4422_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.5 0.255 30.7 ;
      END
   END FE_OFN4422_decrypt

   PIN FE_OFN4476_n_39
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 18 0 18.2 0.255 ;
      END
   END FE_OFN4476_n_39

   PIN FE_OFN4517_n_13659
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.45 0 33.55 0.51 ;
      END
   END FE_OFN4517_n_13659

   PIN FE_OFN4612_n_201
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 3.85 0 3.95 0.51 ;
      END
   END FE_OFN4612_n_201

   PIN FE_OFN4797_n_21953
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 20.55 0.51 20.65 ;
      END
   END FE_OFN4797_n_21953

   PIN FE_OFN663_n_32304
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.85 0 152.95 0.51 ;
      END
   END FE_OFN663_n_32304

   PIN FE_OFN669_n_32833
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.85 0 234.95 0.51 ;
      END
   END FE_OFN669_n_32833

   PIN FE_OFN677_n_30310
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 372.25 0 372.35 0.51 ;
      END
   END FE_OFN677_n_30310

   PIN FE_OFN683_n_117971
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 160.15 0.51 160.25 ;
      END
   END FE_OFN683_n_117971

   PIN FE_OFN692_n_27625
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 171.95 0.51 172.05 ;
      END
   END FE_OFN692_n_27625

   PIN FE_OFN852_n_3353
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 12.25 0 12.35 0.51 ;
      END
   END FE_OFN852_n_3353

   PIN FE_OFN910_n_21872
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 19.95 0.51 20.05 ;
      END
   END FE_OFN910_n_21872

   PIN FE_OFN947_n_3795
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 27.55 0.51 27.65 ;
      END
   END FE_OFN947_n_3795

   PIN FE_OFN972_n_63299
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.15 0.51 16.25 ;
      END
   END FE_OFN972_n_63299

   PIN g205805_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 232.45 0 232.55 0.51 ;
      END
   END g205805_sb

   PIN g231413_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 76.35 0.51 76.45 ;
      END
   END g231413_p

   PIN g233023_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.25 295.49 72.35 296 ;
      END
   END g233023_p

   PIN g233195_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 21.65 0 21.75 0.51 ;
      END
   END g233195_p

   PIN g235329_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.05 0 68.15 0.51 ;
      END
   END g235329_p

   PIN g265215_p2
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 276.25 0 276.35 0.51 ;
      END
   END g265215_p2

   PIN g266100_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.05 0 198.15 0.51 ;
      END
   END g266100_p

   PIN g267780_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 223.65 0 223.75 0.51 ;
      END
   END g267780_p

   PIN g267919_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 236.05 0 236.15 0.51 ;
      END
   END g267919_p

   PIN g268186_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 216.05 0 216.15 0.51 ;
      END
   END g268186_p

   PIN g268308_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 204.65 0 204.75 0.51 ;
      END
   END g268308_p

   PIN g268393_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.65 0 152.75 0.51 ;
      END
   END g268393_p

   PIN g268990_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.65 0 127.75 0.51 ;
      END
   END g268990_p

   PIN g269848_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 358.45 0 358.55 0.51 ;
      END
   END g269848_p

   PIN g270852_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 195.05 0 195.15 0.51 ;
      END
   END g270852_p

   PIN g271549_p1
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 194.45 0 194.55 0.51 ;
      END
   END g271549_p1

   PIN g271686_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.85 0 177.95 0.51 ;
      END
   END g271686_p

   PIN g271749_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 182.45 0 182.55 0.51 ;
      END
   END g271749_p

   PIN g271784_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.05 0 185.15 0.51 ;
      END
   END g271784_p

   PIN g271972_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 195.25 0 195.35 0.51 ;
      END
   END g271972_p

   PIN g272788_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 179.05 0 179.15 0.51 ;
      END
   END g272788_p

   PIN g272818_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 39.85 0 39.95 0.51 ;
      END
   END g272818_sb

   PIN g272848_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.45 0 38.55 0.51 ;
      END
   END g272848_p

   PIN g273938_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 25.95 0.51 26.05 ;
      END
   END g273938_p

   PIN g273953_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.55 0.51 42.65 ;
      END
   END g273953_p

   PIN g278067_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 13.65 0 13.75 0.51 ;
      END
   END g278067_p

   PIN g279539_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.45 0 20.55 0.51 ;
      END
   END g279539_db

   PIN g279539_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.25 0 11.35 0.51 ;
      END
   END g279539_sb

   PIN g302013_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 20.75 0.51 20.85 ;
      END
   END g302013_p

   PIN g302028_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.25 0 3.35 0.51 ;
      END
   END g302028_p

   PIN g302042_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 52.55 0.51 52.65 ;
      END
   END g302042_p

   PIN g302689_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 20.95 0.51 21.05 ;
      END
   END g302689_p

   PIN g303333_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 27.35 0.51 27.45 ;
      END
   END g303333_p

   PIN g303373_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 5.85 0 5.95 0.51 ;
      END
   END g303373_p

   PIN g304261_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.85 0 2.95 0.51 ;
      END
   END g304261_p

   PIN g304290_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 5.65 0 5.75 0.51 ;
      END
   END g304290_p

   PIN g304292_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 7.25 0 7.35 0.51 ;
      END
   END g304292_p

   PIN g305157_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 94.25 0 94.35 0.51 ;
      END
   END g305157_p

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.45 0 41.55 0.51 ;
      END
   END ispd_clk

   PIN key1_19_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.05 295.49 8.15 296 ;
      END
   END key1_19_

   PIN key1_55_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.05 295.49 92.15 296 ;
      END
   END key1_55_

   PIN key3_19_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.05 295.49 12.15 296 ;
      END
   END key3_19_

   PIN key3_55_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.05 295.49 104.15 296 ;
      END
   END key3_55_

   PIN n_1023
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.95 0.51 51.05 ;
      END
   END n_1023

   PIN n_10608
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15.45 0 15.55 0.51 ;
      END
   END n_10608

   PIN n_108553
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.05 0 127.15 0.51 ;
      END
   END n_108553

   PIN n_108562
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 48.15 0.51 48.25 ;
      END
   END n_108562

   PIN n_108697
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.75 0.51 64.85 ;
      END
   END n_108697

   PIN n_108698
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.05 0 92.15 0.51 ;
      END
   END n_108698

   PIN n_108729
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.55 0.51 40.65 ;
      END
   END n_108729

   PIN n_108760
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.25 0 41.35 0.51 ;
      END
   END n_108760

   PIN n_108971
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 14.45 0 14.55 0.51 ;
      END
   END n_108971

   PIN n_109090
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 344.25 0 344.35 0.51 ;
      END
   END n_109090

   PIN n_109137
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.65 0 40.75 0.51 ;
      END
   END n_109137

   PIN n_109138
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.05 0 41.15 0.51 ;
      END
   END n_109138

   PIN n_112756
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.45 295.49 128.55 296 ;
      END
   END n_112756

   PIN n_112757
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.25 295.49 128.35 296 ;
      END
   END n_112757

   PIN n_112829
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.85 0 139.95 0.51 ;
      END
   END n_112829

   PIN n_116914
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 30.45 0 30.55 0.51 ;
      END
   END n_116914

   PIN n_116948
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 51.85 0 51.95 0.51 ;
      END
   END n_116948

   PIN n_117298
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.05 0 166.15 0.51 ;
      END
   END n_117298

   PIN n_117339
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.25 0 18.35 0.51 ;
      END
   END n_117339

   PIN n_117340
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 52.75 0.51 52.85 ;
      END
   END n_117340

   PIN n_117465
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 40.05 0 40.15 0.51 ;
      END
   END n_117465

   PIN n_117466
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 21.45 0 21.55 0.51 ;
      END
   END n_117466

   PIN n_117596
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 224.25 0 224.35 0.51 ;
      END
   END n_117596

   PIN n_117600
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 207.65 0 207.75 0.51 ;
      END
   END n_117600

   PIN n_117902
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.35 0.51 28.45 ;
      END
   END n_117902

   PIN n_118304
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 143.25 0 143.35 0.51 ;
      END
   END n_118304

   PIN n_118305
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 142.65 0 142.75 0.51 ;
      END
   END n_118305

   PIN n_118591
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 16.65 295.49 16.75 296 ;
      END
   END n_118591

   PIN n_118596
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.45 0 8.55 0.51 ;
      END
   END n_118596

   PIN n_118598
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 18.05 295.49 18.15 296 ;
      END
   END n_118598

   PIN n_1263
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 16.45 0 16.55 0.51 ;
      END
   END n_1263

   PIN n_1266
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 13.45 0 13.55 0.51 ;
      END
   END n_1266

   PIN n_1281
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.95 0.51 16.05 ;
      END
   END n_1281

   PIN n_1387
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.45 0 28.55 0.51 ;
      END
   END n_1387

   PIN n_13938
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.65 0 15.75 0.51 ;
      END
   END n_13938

   PIN n_1489
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 50.95 0.51 51.05 ;
      END
   END n_1489

   PIN n_1501
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.45 0 15.55 0.51 ;
      END
   END n_1501

   PIN n_1504
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 12.25 0 12.35 0.51 ;
      END
   END n_1504

   PIN n_1529
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 5.45 0 5.55 0.51 ;
      END
   END n_1529

   PIN n_155186
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.85 0 127.95 0.51 ;
      END
   END n_155186

   PIN n_1593
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.95 0.51 34.05 ;
      END
   END n_1593

   PIN n_1646
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 11.15 0.51 11.25 ;
      END
   END n_1646

   PIN n_18158
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.35 0.51 22.45 ;
      END
   END n_18158

   PIN n_18380
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 3.05 0 3.15 0.51 ;
      END
   END n_18380

   PIN n_18386
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.35 0.51 31.45 ;
      END
   END n_18386

   PIN n_1848
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 24.65 0 24.75 0.51 ;
      END
   END n_1848

   PIN n_18639
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 12.05 0 12.15 0.51 ;
      END
   END n_18639

   PIN n_18670
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.65 0 21.75 0.51 ;
      END
   END n_18670

   PIN n_18679
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 219.95 0.51 220.05 ;
      END
   END n_18679

   PIN n_1878
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.25 0 6.35 0.51 ;
      END
   END n_1878

   PIN n_18862
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.15 0.51 21.25 ;
      END
   END n_18862

   PIN n_19056
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 2.85 0 2.95 0.51 ;
      END
   END n_19056

   PIN n_19424
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.65 0 4.75 0.51 ;
      END
   END n_19424

   PIN n_19436
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.15 0.51 35.25 ;
      END
   END n_19436

   PIN n_19692
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.35 0.51 27.45 ;
      END
   END n_19692

   PIN n_19693
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.75 0.51 15.85 ;
      END
   END n_19693

   PIN n_19844
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 208.15 0.51 208.25 ;
      END
   END n_19844

   PIN n_19868
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.05 0 6.15 0.51 ;
      END
   END n_19868

   PIN n_20239
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 29.15 0.51 29.25 ;
      END
   END n_20239

   PIN n_20284
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 207.95 0.51 208.05 ;
      END
   END n_20284

   PIN n_20529
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.55 0.51 15.65 ;
      END
   END n_20529

   PIN n_20542
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.35 0.51 15.45 ;
      END
   END n_20542

   PIN n_20744
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.45 0 4.55 0.51 ;
      END
   END n_20744

   PIN n_20818
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 20.15 0.51 20.25 ;
      END
   END n_20818

   PIN n_21311
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.45 0 14.55 0.51 ;
      END
   END n_21311

   PIN n_2155
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.05 0 5.15 0.51 ;
      END
   END n_2155

   PIN n_21823
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.15 0.51 36.25 ;
      END
   END n_21823

   PIN n_21905
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.35 0.51 21.45 ;
      END
   END n_21905

   PIN n_21912
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.45 0 26.55 0.51 ;
      END
   END n_21912

   PIN n_21921
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 243.55 0.51 243.65 ;
      END
   END n_21921

   PIN n_21949
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.35 0.51 62.45 ;
      END
   END n_21949

   PIN n_21999
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.05 0 22.15 0.51 ;
      END
   END n_21999

   PIN n_22036
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.15 0.51 51.25 ;
      END
   END n_22036

   PIN n_22173
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 24.25 0 24.35 0.51 ;
      END
   END n_22173

   PIN n_22174
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.25 0 20.35 0.51 ;
      END
   END n_22174

   PIN n_22255
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.25 0 20.35 0.51 ;
      END
   END n_22255

   PIN n_22325
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 24.45 0 24.55 0.51 ;
      END
   END n_22325

   PIN n_22338
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 41.25 0 41.35 0.51 ;
      END
   END n_22338

   PIN n_22350
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.85 0 17.95 0.51 ;
      END
   END n_22350

   PIN n_22352
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 16.05 0 16.15 0.51 ;
      END
   END n_22352

   PIN n_22359
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.25 0 22.35 0.51 ;
      END
   END n_22359

   PIN n_22392
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 1.85 0 1.95 0.51 ;
      END
   END n_22392

   PIN n_22454
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 52.95 0.51 53.05 ;
      END
   END n_22454

   PIN n_22603
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.15 0.51 30.25 ;
      END
   END n_22603

   PIN n_22612
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 30.95 0.51 31.05 ;
      END
   END n_22612

   PIN n_22800
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 15.05 0 15.15 0.51 ;
      END
   END n_22800

   PIN n_22836
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 40.35 0.51 40.45 ;
      END
   END n_22836

   PIN n_22929
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 40.55 0.51 40.65 ;
      END
   END n_22929

   PIN n_22932
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 19.25 0 19.35 0.51 ;
      END
   END n_22932

   PIN n_22937
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 36.55 0.51 36.65 ;
      END
   END n_22937

   PIN n_23053
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.65 0 23.75 0.51 ;
      END
   END n_23053

   PIN n_23062
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 14.25 0 14.35 0.51 ;
      END
   END n_23062

   PIN n_23073
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.65 0 19.75 0.51 ;
      END
   END n_23073

   PIN n_23091
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.85 0 20.95 0.51 ;
      END
   END n_23091

   PIN n_23165
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 53.15 0.51 53.25 ;
      END
   END n_23165

   PIN n_23219
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 26.75 0.51 26.85 ;
      END
   END n_23219

   PIN n_2332
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 21.05 0 21.15 0.51 ;
      END
   END n_2332

   PIN n_2334
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.95 0.51 65.05 ;
      END
   END n_2334

   PIN n_23606
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.65 0 22.75 0.51 ;
      END
   END n_23606

   PIN n_23635
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 19.65 0 19.75 0.51 ;
      END
   END n_23635

   PIN n_23694
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.05 0 27.15 0.51 ;
      END
   END n_23694

   PIN n_23721
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 26.85 0 26.95 0.51 ;
      END
   END n_23721

   PIN n_23876
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.55 0.51 21.65 ;
      END
   END n_23876

   PIN n_24030
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.75 0.51 21.85 ;
      END
   END n_24030

   PIN n_24048
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 10.75 0.51 10.85 ;
      END
   END n_24048

   PIN n_2435
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.15 0.51 15.25 ;
      END
   END n_2435

   PIN n_24781
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.95 0.51 15.05 ;
      END
   END n_24781

   PIN n_2483
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.45 0 16.55 0.51 ;
      END
   END n_2483

   PIN n_2504
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 6.45 0 6.55 0.51 ;
      END
   END n_2504

   PIN n_25070
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 13.15 0.51 13.25 ;
      END
   END n_25070

   PIN n_25088
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.25 295.49 56.35 296 ;
      END
   END n_25088

   PIN n_25090
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44.05 295.49 44.15 296 ;
      END
   END n_25090

   PIN n_25102
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.65 295.49 3.75 296 ;
      END
   END n_25102

   PIN n_25130
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 2.65 295.49 2.75 296 ;
      END
   END n_25130

   PIN n_25224
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.55 0.51 23.65 ;
      END
   END n_25224

   PIN n_25227
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.75 0.51 14.85 ;
      END
   END n_25227

   PIN n_25228
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.15 0.51 28.25 ;
      END
   END n_25228

   PIN n_25317
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.35 0.51 23.45 ;
      END
   END n_25317

   PIN n_25375
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.55 0.51 14.65 ;
      END
   END n_25375

   PIN n_25412
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.15 0.51 23.25 ;
      END
   END n_25412

   PIN n_2549
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 39.65 0 39.75 0.51 ;
      END
   END n_2549

   PIN n_25591
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.25 295.49 44.35 296 ;
      END
   END n_25591

   PIN n_25662
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 62.95 0.51 63.05 ;
      END
   END n_25662

   PIN n_25669
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.05 295.49 44.15 296 ;
      END
   END n_25669

   PIN n_25671
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.85 295.49 55.95 296 ;
      END
   END n_25671

   PIN n_25677
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.85 295.49 43.95 296 ;
      END
   END n_25677

   PIN n_25679
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.85 295.49 16.95 296 ;
      END
   END n_25679

   PIN n_25713
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.85 295.49 55.95 296 ;
      END
   END n_25713

   PIN n_25727
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 75.75 0.51 75.85 ;
      END
   END n_25727

   PIN n_25764
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 76.15 0.51 76.25 ;
      END
   END n_25764

   PIN n_25771
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 12.75 0.51 12.85 ;
      END
   END n_25771

   PIN n_25794
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.25 0 6.35 0.51 ;
      END
   END n_25794

   PIN n_25810
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 114.85 0 114.95 0.51 ;
      END
   END n_25810

   PIN n_25823
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.35 0.51 44.45 ;
      END
   END n_25823

   PIN n_25837
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 90.65 0 90.75 0.51 ;
      END
   END n_25837

   PIN n_25849
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.05 0 38.15 0.51 ;
      END
   END n_25849

   PIN n_25856
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 19.85 0 19.95 0.51 ;
      END
   END n_25856

   PIN n_25870
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 25.85 0 25.95 0.51 ;
      END
   END n_25870

   PIN n_25888
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 32.25 0 32.35 0.51 ;
      END
   END n_25888

   PIN n_25889
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.15 0.51 25.25 ;
      END
   END n_25889

   PIN n_25895
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 26.55 0.51 26.65 ;
      END
   END n_25895

   PIN n_25935
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 186.25 0 186.35 0.51 ;
      END
   END n_25935

   PIN n_26069
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 46.85 0 46.95 0.51 ;
      END
   END n_26069

   PIN n_26071
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.55 0.51 44.65 ;
      END
   END n_26071

   PIN n_26153
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.05 295.49 80.15 296 ;
      END
   END n_26153

   PIN n_26374
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 24.75 0.51 24.85 ;
      END
   END n_26374

   PIN n_26377
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.75 0.51 9.85 ;
      END
   END n_26377

   PIN n_26491
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.25 0 91.35 0.51 ;
      END
   END n_26491

   PIN n_26510
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.45 0 55.55 0.51 ;
      END
   END n_26510

   PIN n_26547
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.9 0.255 43.1 ;
      END
   END n_26547

   PIN n_26553
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.35 0.51 50.45 ;
      END
   END n_26553

   PIN n_26558
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 7.05 0 7.15 0.51 ;
      END
   END n_26558

   PIN n_26622
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 47.95 0.51 48.05 ;
      END
   END n_26622

   PIN n_2663
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 78.65 0 78.75 0.51 ;
      END
   END n_2663

   PIN n_26632
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 41.75 0.51 41.85 ;
      END
   END n_26632

   PIN n_26638
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 8.95 0.51 9.05 ;
      END
   END n_26638

   PIN n_26672
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 45.15 0.51 45.25 ;
      END
   END n_26672

   PIN n_26763
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.95 0.51 44.05 ;
      END
   END n_26763

   PIN n_26765
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 44.95 0.51 45.05 ;
      END
   END n_26765

   PIN n_26785
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.55 0.51 43.65 ;
      END
   END n_26785

   PIN n_2679
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 13.55 0.51 13.65 ;
      END
   END n_2679

   PIN n_26983
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.75 0.51 40.85 ;
      END
   END n_26983

   PIN n_27075
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.15 0.51 42.25 ;
      END
   END n_27075

   PIN n_2708
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 26.95 0.51 27.05 ;
      END
   END n_2708

   PIN n_27099
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 4.05 0 4.15 0.51 ;
      END
   END n_27099

   PIN n_27127
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 9.15 0.51 9.25 ;
      END
   END n_27127

   PIN n_27563
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 21.55 0.51 21.65 ;
      END
   END n_27563

   PIN n_27603
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.55 0.51 87.65 ;
      END
   END n_27603

   PIN n_27616
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.85 0 24.95 0.51 ;
      END
   END n_27616

   PIN n_27646
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 63.75 0.51 63.85 ;
      END
   END n_27646

   PIN n_27654
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 90.45 0 90.55 0.51 ;
      END
   END n_27654

   PIN n_27671
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 232.15 0.51 232.25 ;
      END
   END n_27671

   PIN n_27702
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 220.15 0.51 220.25 ;
      END
   END n_27702

   PIN n_27743
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 38.75 0.51 38.85 ;
      END
   END n_27743

   PIN n_27794
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.25 0 36.35 0.51 ;
      END
   END n_27794

   PIN n_2780
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.35 0.51 14.45 ;
      END
   END n_2780

   PIN n_27806
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 36.05 0 36.15 0.51 ;
      END
   END n_27806

   PIN n_27815
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 58.85 0 58.95 0.51 ;
      END
   END n_27815

   PIN n_27847
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 18.85 0 18.95 0.51 ;
      END
   END n_27847

   PIN n_27858
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.45 0 319.55 0.51 ;
      END
   END n_27858

   PIN n_27869
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 260.05 0 260.15 0.51 ;
      END
   END n_27869

   PIN n_27978
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.25 0 103.35 0.51 ;
      END
   END n_27978

   PIN n_27984
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.65 0 103.75 0.51 ;
      END
   END n_27984

   PIN n_28031
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.25 0 101.35 0.51 ;
      END
   END n_28031

   PIN n_28036
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 105.25 0 105.35 0.51 ;
      END
   END n_28036

   PIN n_28044
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 99.45 0 99.55 0.51 ;
      END
   END n_28044

   PIN n_28072
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.25 0 102.35 0.51 ;
      END
   END n_28072

   PIN n_281
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 10.95 0.51 11.05 ;
      END
   END n_281

   PIN n_28101
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.05 0 115.15 0.51 ;
      END
   END n_28101

   PIN n_28135
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.25 0 164.35 0.51 ;
      END
   END n_28135

   PIN n_28136
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.65 0 163.75 0.51 ;
      END
   END n_28136

   PIN n_28138
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 177.85 0 177.95 0.51 ;
      END
   END n_28138

   PIN n_28140
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 180.45 0 180.55 0.51 ;
      END
   END n_28140

   PIN n_28166
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 39.85 0 39.95 0.51 ;
      END
   END n_28166

   PIN n_28204
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.05 0 175.15 0.51 ;
      END
   END n_28204

   PIN n_28212
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 92.65 0 92.75 0.51 ;
      END
   END n_28212

   PIN n_28230
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 107.25 0 107.35 0.51 ;
      END
   END n_28230

   PIN n_28237
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 102.8 0 103 0.255 ;
      END
   END n_28237

   PIN n_28309
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 102.4 0 102.6 0.255 ;
      END
   END n_28309

   PIN n_28396
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 190.65 0 190.75 0.51 ;
      END
   END n_28396

   PIN n_28398
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 105.45 0 105.55 0.51 ;
      END
   END n_28398

   PIN n_28447
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.85 0 103.95 0.51 ;
      END
   END n_28447

   PIN n_28448
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 183.65 0 183.75 0.51 ;
      END
   END n_28448

   PIN n_28501
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.05 0 116.15 0.51 ;
      END
   END n_28501

   PIN n_28504
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 101.85 0 101.95 0.51 ;
      END
   END n_28504

   PIN n_28534
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.45 0 115.55 0.51 ;
      END
   END n_28534

   PIN n_28606
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 102.05 0 102.15 0.51 ;
      END
   END n_28606

   PIN n_28621
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.85 0 114.95 0.51 ;
      END
   END n_28621

   PIN n_28622
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 96.25 0 96.35 0.51 ;
      END
   END n_28622

   PIN n_28639
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 183.45 0 183.55 0.51 ;
      END
   END n_28639

   PIN n_28712
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.25 0 104.35 0.51 ;
      END
   END n_28712

   PIN n_28713
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.45 0 100.55 0.51 ;
      END
   END n_28713

   PIN n_28715
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 99.25 0 99.35 0.51 ;
      END
   END n_28715

   PIN n_28717
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.05 0 98.15 0.51 ;
      END
   END n_28717

   PIN n_28780
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.85 0 115.95 0.51 ;
      END
   END n_28780

   PIN n_28805
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 114.65 0 114.75 0.51 ;
      END
   END n_28805

   PIN n_28859
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.85 0 102.95 0.51 ;
      END
   END n_28859

   PIN n_2887
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 62.75 0.51 62.85 ;
      END
   END n_2887

   PIN n_28880
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 193.05 0 193.15 0.51 ;
      END
   END n_28880

   PIN n_29030
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 187.45 0 187.55 0.51 ;
      END
   END n_29030

   PIN n_29061
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.85 0 93.95 0.51 ;
      END
   END n_29061

   PIN n_29110
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.85 0 176.95 0.51 ;
      END
   END n_29110

   PIN n_29123
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 98.85 0 98.95 0.51 ;
      END
   END n_29123

   PIN n_29127
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 114.25 0 114.35 0.51 ;
      END
   END n_29127

   PIN n_29141
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 182.25 0 182.35 0.51 ;
      END
   END n_29141

   PIN n_29150
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 195.05 0 195.15 0.51 ;
      END
   END n_29150

   PIN n_29151
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.85 0 185.95 0.51 ;
      END
   END n_29151

   PIN n_29239
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 103.85 0 103.95 0.51 ;
      END
   END n_29239

   PIN n_29241
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 183.85 0 183.95 0.51 ;
      END
   END n_29241

   PIN n_29246
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 185.85 0 185.95 0.51 ;
      END
   END n_29246

   PIN n_29249
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 182.85 0 182.95 0.51 ;
      END
   END n_29249

   PIN n_29264
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.85 0 188.95 0.51 ;
      END
   END n_29264

   PIN n_29280
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 186.45 0 186.55 0.51 ;
      END
   END n_29280

   PIN n_29332
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 178.25 0 178.35 0.51 ;
      END
   END n_29332

   PIN n_29350
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 181.85 0 181.95 0.51 ;
      END
   END n_29350

   PIN n_29362
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 102.45 0 102.55 0.51 ;
      END
   END n_29362

   PIN n_29371
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 183.05 0 183.15 0.51 ;
      END
   END n_29371

   PIN n_29378
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 179.45 0 179.55 0.51 ;
      END
   END n_29378

   PIN n_29461
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.45 0 177.55 0.51 ;
      END
   END n_29461

   PIN n_29470
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.65 0 171.75 0.51 ;
      END
   END n_29470

   PIN n_29524
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 115.25 0 115.35 0.51 ;
      END
   END n_29524

   PIN n_29539
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.05 0 104.15 0.51 ;
      END
   END n_29539

   PIN n_29544
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 180.05 0 180.15 0.51 ;
      END
   END n_29544

   PIN n_29549
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 171.45 0 171.55 0.51 ;
      END
   END n_29549

   PIN n_29562
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 103.45 0 103.55 0.51 ;
      END
   END n_29562

   PIN n_29593
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 101.85 0 101.95 0.51 ;
      END
   END n_29593

   PIN n_29594
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 77.65 0 77.75 0.51 ;
      END
   END n_29594

   PIN n_29595
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 101.65 0 101.75 0.51 ;
      END
   END n_29595

   PIN n_29611
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 93.05 0 93.15 0.51 ;
      END
   END n_29611

   PIN n_29645
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 77.05 0 77.15 0.51 ;
      END
   END n_29645

   PIN n_29649
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.05 0 93.15 0.51 ;
      END
   END n_29649

   PIN n_29753
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 198.65 0 198.75 0.51 ;
      END
   END n_29753

   PIN n_29756
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 103.25 0 103.35 0.51 ;
      END
   END n_29756

   PIN n_29817
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 127.25 0 127.35 0.51 ;
      END
   END n_29817

   PIN n_29840
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 295.65 0 295.75 0.51 ;
      END
   END n_29840

   PIN n_29877
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 379.25 0 379.35 0.51 ;
      END
   END n_29877

   PIN n_29906
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 339.65 0 339.75 0.51 ;
      END
   END n_29906

   PIN n_29918
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 113.45 0 113.55 0.51 ;
      END
   END n_29918

   PIN n_29943
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 175.85 0 175.95 0.51 ;
      END
   END n_29943

   PIN n_29949
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 335.45 0 335.55 0.51 ;
      END
   END n_29949

   PIN n_29998
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 392.25 0 392.35 0.51 ;
      END
   END n_29998

   PIN n_30001
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 335.05 0 335.15 0.51 ;
      END
   END n_30001

   PIN n_30010
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 121.85 0 121.95 0.51 ;
      END
   END n_30010

   PIN n_30013
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 333.45 0 333.55 0.51 ;
      END
   END n_30013

   PIN n_30018
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 114.45 0 114.55 0.51 ;
      END
   END n_30018

   PIN n_30045
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 343.05 0 343.15 0.51 ;
      END
   END n_30045

   PIN n_30049
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 404.05 0 404.15 0.51 ;
      END
   END n_30049

   PIN n_30051
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 380.05 0 380.15 0.51 ;
      END
   END n_30051

   PIN n_30107
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 371.45 0 371.55 0.51 ;
      END
   END n_30107

   PIN n_30111
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.05 0 139.15 0.51 ;
      END
   END n_30111

   PIN n_30142
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.2 0 163.4 0.255 ;
      END
   END n_30142

   PIN n_30206
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 329.25 0 329.35 0.51 ;
      END
   END n_30206

   PIN n_30225
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 138.85 0 138.95 0.51 ;
      END
   END n_30225

   PIN n_30242
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 363.85 0 363.95 0.51 ;
      END
   END n_30242

   PIN n_30259
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 379.45 0 379.55 0.51 ;
      END
   END n_30259

   PIN n_30263
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 415.85 0 415.95 0.51 ;
      END
   END n_30263

   PIN n_30295
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 366.65 0 366.75 0.51 ;
      END
   END n_30295

   PIN n_30358
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 326.85 0 326.95 0.51 ;
      END
   END n_30358

   PIN n_30390
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 374.85 0 374.95 0.51 ;
      END
   END n_30390

   PIN n_30400
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 355.45 0 355.55 0.51 ;
      END
   END n_30400

   PIN n_30406
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 355.25 0 355.35 0.51 ;
      END
   END n_30406

   PIN n_30418
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 379.45 0 379.55 0.51 ;
      END
   END n_30418

   PIN n_3045
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 14.65 0 14.75 0.51 ;
      END
   END n_3045

   PIN n_30454
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 338.25 0 338.35 0.51 ;
      END
   END n_30454

   PIN n_30461
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 333.05 0 333.15 0.51 ;
      END
   END n_30461

   PIN n_30527
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 372.05 0 372.15 0.51 ;
      END
   END n_30527

   PIN n_30528
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 360.25 0 360.35 0.51 ;
      END
   END n_30528

   PIN n_30544
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 379.65 0 379.75 0.51 ;
      END
   END n_30544

   PIN n_30655
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 334.45 0 334.55 0.51 ;
      END
   END n_30655

   PIN n_30686
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 392.45 0 392.55 0.51 ;
      END
   END n_30686

   PIN n_30726
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 365.65 0 365.75 0.51 ;
      END
   END n_30726

   PIN n_30745
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 432.25 0 432.35 0.51 ;
      END
   END n_30745

   PIN n_30755
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 355.05 0 355.15 0.51 ;
      END
   END n_30755

   PIN n_30780
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 379.65 0 379.75 0.51 ;
      END
   END n_30780

   PIN n_30792
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 380.25 0 380.35 0.51 ;
      END
   END n_30792

   PIN n_30818
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 126.8 0 127 0.255 ;
      END
   END n_30818

   PIN n_30835
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 416.05 0 416.15 0.51 ;
      END
   END n_30835

   PIN n_30917
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 341.65 0 341.75 0.51 ;
      END
   END n_30917

   PIN n_30997
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 376.05 0 376.15 0.51 ;
      END
   END n_30997

   PIN n_31021
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 380.45 0 380.55 0.51 ;
      END
   END n_31021

   PIN n_31023
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 359.85 0 359.95 0.51 ;
      END
   END n_31023

   PIN n_31039
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 392.25 0 392.35 0.51 ;
      END
   END n_31039

   PIN n_31077
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 332.85 0 332.95 0.51 ;
      END
   END n_31077

   PIN n_31091
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 344.45 0 344.55 0.51 ;
      END
   END n_31091

   PIN n_31095
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 357.65 0 357.75 0.51 ;
      END
   END n_31095

   PIN n_31106
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.65 0 140.75 0.51 ;
      END
   END n_31106

   PIN n_31114
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 126.45 0 126.55 0.51 ;
      END
   END n_31114

   PIN n_31122
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 392.65 0 392.75 0.51 ;
      END
   END n_31122

   PIN n_31130
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 146.25 0 146.35 0.51 ;
      END
   END n_31130

   PIN n_31132
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 356.65 0 356.75 0.51 ;
      END
   END n_31132

   PIN n_31146
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 339.65 0 339.75 0.51 ;
      END
   END n_31146

   PIN n_31149
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 342.45 0 342.55 0.51 ;
      END
   END n_31149

   PIN n_31165
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.65 0 139.75 0.51 ;
      END
   END n_31165

   PIN n_31179
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.45 0 127.55 0.51 ;
      END
   END n_31179

   PIN n_31222
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 404.05 0 404.15 0.51 ;
      END
   END n_31222

   PIN n_31280
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 342.85 0 342.95 0.51 ;
      END
   END n_31280

   PIN n_31288
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 174.25 0 174.35 0.51 ;
      END
   END n_31288

   PIN n_31304
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 339.85 0 339.95 0.51 ;
      END
   END n_31304

   PIN n_31306
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 341.05 0 341.15 0.51 ;
      END
   END n_31306

   PIN n_31333
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 145.85 0 145.95 0.51 ;
      END
   END n_31333

   PIN n_31342
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 132.25 0 132.35 0.51 ;
      END
   END n_31342

   PIN n_31345
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.45 0 126.55 0.51 ;
      END
   END n_31345

   PIN n_3136
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 63.95 0.51 64.05 ;
      END
   END n_3136

   PIN n_31381
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 132.05 0 132.15 0.51 ;
      END
   END n_31381

   PIN n_31430
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.05 0 151.15 0.51 ;
      END
   END n_31430

   PIN n_31463
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.25 0 127.35 0.51 ;
      END
   END n_31463

   PIN n_31464
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 329.05 0 329.15 0.51 ;
      END
   END n_31464

   PIN n_31479
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.85 0 139.95 0.51 ;
      END
   END n_31479

   PIN n_31497
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 324.45 0 324.55 0.51 ;
      END
   END n_31497

   PIN n_31510
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 354.25 0 354.35 0.51 ;
      END
   END n_31510

   PIN n_31514
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 144.05 0 144.15 0.51 ;
      END
   END n_31514

   PIN n_31533
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.65 0 115.75 0.51 ;
      END
   END n_31533

   PIN n_31543
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 359.25 0 359.35 0.51 ;
      END
   END n_31543

   PIN n_31544
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 359.05 0 359.15 0.51 ;
      END
   END n_31544

   PIN n_31547
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 355.85 0 355.95 0.51 ;
      END
   END n_31547

   PIN n_31552
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 344.05 0 344.15 0.51 ;
      END
   END n_31552

   PIN n_31587
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.25 0 126.35 0.51 ;
      END
   END n_31587

   PIN n_31609
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.05 0 126.15 0.51 ;
      END
   END n_31609

   PIN n_31644
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 152.25 0 152.35 0.51 ;
      END
   END n_31644

   PIN n_3165
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.55 0.51 12.65 ;
      END
   END n_3165

   PIN n_31657
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 345.45 0 345.55 0.51 ;
      END
   END n_31657

   PIN n_31659
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.65 0 139.75 0.51 ;
      END
   END n_31659

   PIN n_31667
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 125.85 0 125.95 0.51 ;
      END
   END n_31667

   PIN n_31668
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.05 0 139.15 0.51 ;
      END
   END n_31668

   PIN n_31669
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.85 0 138.95 0.51 ;
      END
   END n_31669

   PIN n_31684
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 345.25 0 345.35 0.51 ;
      END
   END n_31684

   PIN n_31685
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 233.85 0 233.95 0.51 ;
      END
   END n_31685

   PIN n_31701
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.85 0 308.95 0.51 ;
      END
   END n_31701

   PIN n_31716
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 313.25 0 313.35 0.51 ;
      END
   END n_31716

   PIN n_31733
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.25 0 139.35 0.51 ;
      END
   END n_31733

   PIN n_31742
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.85 0 267.95 0.51 ;
      END
   END n_31742

   PIN n_31745
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 260.25 0 260.35 0.51 ;
      END
   END n_31745

   PIN n_31829
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 160.85 0 160.95 0.51 ;
      END
   END n_31829

   PIN n_31855
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 216.85 0 216.95 0.51 ;
      END
   END n_31855

   PIN n_31857
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 222.85 0 222.95 0.51 ;
      END
   END n_31857

   PIN n_3189
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 26.35 0.51 26.45 ;
      END
   END n_3189

   PIN n_31896
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 162.65 0 162.75 0.51 ;
      END
   END n_31896

   PIN n_31898
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 214.05 0 214.15 0.51 ;
      END
   END n_31898

   PIN n_31911
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 201.05 0 201.15 0.51 ;
      END
   END n_31911

   PIN n_32023
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 312.25 0 312.35 0.51 ;
      END
   END n_32023

   PIN n_32055
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 247.85 0 247.95 0.51 ;
      END
   END n_32055

   PIN n_32071
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 207.45 0 207.55 0.51 ;
      END
   END n_32071

   PIN n_32181
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 172.45 0 172.55 0.51 ;
      END
   END n_32181

   PIN n_32200
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 213.65 0 213.75 0.51 ;
      END
   END n_32200

   PIN n_32218
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 259.65 0 259.75 0.51 ;
      END
   END n_32218

   PIN n_32268
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.25 0 212.35 0.51 ;
      END
   END n_32268

   PIN n_32272
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 200.05 0 200.15 0.51 ;
      END
   END n_32272

   PIN n_32333
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 203.25 0 203.35 0.51 ;
      END
   END n_32333

   PIN n_32511
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 215.85 0 215.95 0.51 ;
      END
   END n_32511

   PIN n_32526
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.65 0 132.75 0.51 ;
      END
   END n_32526

   PIN n_32586
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 207.65 0 207.75 0.51 ;
      END
   END n_32586

   PIN n_32608
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.05 0 136.15 0.51 ;
      END
   END n_32608

   PIN n_32620
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 202.85 0 202.95 0.51 ;
      END
   END n_32620

   PIN n_32650
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.25 0 224.35 0.51 ;
      END
   END n_32650

   PIN n_32654
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 218.45 0 218.55 0.51 ;
      END
   END n_32654

   PIN n_32662
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 203.05 0 203.15 0.51 ;
      END
   END n_32662

   PIN n_32677
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 203.05 0 203.15 0.51 ;
      END
   END n_32677

   PIN n_32678
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 259.65 0 259.75 0.51 ;
      END
   END n_32678

   PIN n_32695
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.85 0 224.95 0.51 ;
      END
   END n_32695

   PIN n_32766
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 225.05 0 225.15 0.51 ;
      END
   END n_32766

   PIN n_32777
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.45 0 151.55 0.51 ;
      END
   END n_32777

   PIN n_32803
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 217.65 0 217.75 0.51 ;
      END
   END n_32803

   PIN n_32804
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 226.65 0 226.75 0.51 ;
      END
   END n_32804

   PIN n_32807
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 222.25 0 222.35 0.51 ;
      END
   END n_32807

   PIN n_32810
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 199.65 0 199.75 0.51 ;
      END
   END n_32810

   PIN n_32811
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.45 0 152.55 0.51 ;
      END
   END n_32811

   PIN n_32828
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 207.45 0 207.55 0.51 ;
      END
   END n_32828

   PIN n_32865
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 207.25 0 207.35 0.51 ;
      END
   END n_32865

   PIN n_32866
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 318.6 0 318.8 0.255 ;
      END
   END n_32866

   PIN n_32927
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 206.85 0 206.95 0.51 ;
      END
   END n_32927

   PIN n_32952
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 215.45 0 215.55 0.51 ;
      END
   END n_32952

   PIN n_32970
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.85 0 197.95 0.51 ;
      END
   END n_32970

   PIN n_32976
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 198.05 0 198.15 0.51 ;
      END
   END n_32976

   PIN n_33002
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 235.65 0 235.75 0.51 ;
      END
   END n_33002

   PIN n_33019
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 201.05 0 201.15 0.51 ;
      END
   END n_33019

   PIN n_33073
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 219.45 0 219.55 0.51 ;
      END
   END n_33073

   PIN n_33080
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 227.25 0 227.35 0.51 ;
      END
   END n_33080

   PIN n_33098
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 219.65 0 219.75 0.51 ;
      END
   END n_33098

   PIN n_33134
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 209.05 0 209.15 0.51 ;
      END
   END n_33134

   PIN n_33154
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 198.25 0 198.35 0.51 ;
      END
   END n_33154

   PIN n_33172
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.25 0 152.35 0.51 ;
      END
   END n_33172

   PIN n_33210
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.05 0 220.15 0.51 ;
      END
   END n_33210

   PIN n_33229
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.25 0 211.35 0.51 ;
      END
   END n_33229

   PIN n_33295
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 222.05 0 222.15 0.51 ;
      END
   END n_33295

   PIN n_33371
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 208.65 0 208.75 0.51 ;
      END
   END n_33371

   PIN n_33389
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.05 0 152.15 0.51 ;
      END
   END n_33389

   PIN n_33406
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.45 0 132.55 0.51 ;
      END
   END n_33406

   PIN n_33437
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.65 0 136.75 0.51 ;
      END
   END n_33437

   PIN n_33472
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.85 0 136.95 0.51 ;
      END
   END n_33472

   PIN n_33499
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 134.05 0 134.15 0.51 ;
      END
   END n_33499

   PIN n_3351
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.75 0.51 31.85 ;
      END
   END n_3351

   PIN n_33543
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 199.05 0 199.15 0.51 ;
      END
   END n_33543

   PIN n_33601
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.85 0 124.95 0.51 ;
      END
   END n_33601

   PIN n_33602
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.45 0 139.55 0.51 ;
      END
   END n_33602

   PIN n_33603
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.45 0 139.55 0.51 ;
      END
   END n_33603

   PIN n_33604
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.25 0 139.35 0.51 ;
      END
   END n_33604

   PIN n_33627
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 252.05 0 252.15 0.51 ;
      END
   END n_33627

   PIN n_33638
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 198.45 0 198.55 0.51 ;
      END
   END n_33638

   PIN n_33667
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 197.85 0 197.95 0.51 ;
      END
   END n_33667

   PIN n_33701
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.65 0 197.75 0.51 ;
      END
   END n_33701

   PIN n_33735
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.45 0 163.55 0.51 ;
      END
   END n_33735

   PIN n_33977
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.05 0 272.15 0.51 ;
      END
   END n_33977

   PIN n_34040
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 288.85 0 288.95 0.51 ;
      END
   END n_34040

   PIN n_34127
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.65 0 285.75 0.51 ;
      END
   END n_34127

   PIN n_34204
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.45 0 282.55 0.51 ;
      END
   END n_34204

   PIN n_34217
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 297.25 0 297.35 0.51 ;
      END
   END n_34217

   PIN n_34298
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.25 0 260.35 0.51 ;
      END
   END n_34298

   PIN n_34312
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 280.25 0 280.35 0.51 ;
      END
   END n_34312

   PIN n_34315
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.05 0 285.15 0.51 ;
      END
   END n_34315

   PIN n_34369
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.65 0 272.75 0.51 ;
      END
   END n_34369

   PIN n_34418
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.05 0 293.15 0.51 ;
      END
   END n_34418

   PIN n_34420
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.25 0 281.35 0.51 ;
      END
   END n_34420

   PIN n_34475
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 287.85 0 287.95 0.51 ;
      END
   END n_34475

   PIN n_34501
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.25 0 271.35 0.51 ;
      END
   END n_34501

   PIN n_34505
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 282.2 0 282.4 0.255 ;
      END
   END n_34505

   PIN n_3452
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.95 0.51 33.05 ;
      END
   END n_3452

   PIN n_34605
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 283.05 0 283.15 0.51 ;
      END
   END n_34605

   PIN n_34738
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.85 0 270.95 0.51 ;
      END
   END n_34738

   PIN n_34794
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 286.25 0 286.35 0.51 ;
      END
   END n_34794

   PIN n_34839
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 297.65 0 297.75 0.51 ;
      END
   END n_34839

   PIN n_34903
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 295.65 0 295.75 0.51 ;
      END
   END n_34903

   PIN n_34918
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 297.05 0 297.15 0.51 ;
      END
   END n_34918

   PIN n_34999
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 288.05 0 288.15 0.51 ;
      END
   END n_34999

   PIN n_35106
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 296.65 0 296.75 0.51 ;
      END
   END n_35106

   PIN n_35141
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.25 0 284.35 0.51 ;
      END
   END n_35141

   PIN n_35319
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 278.05 0 278.15 0.51 ;
      END
   END n_35319

   PIN n_3533
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.35 0.51 75.45 ;
      END
   END n_3533

   PIN n_35567
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 299.45 0 299.55 0.51 ;
      END
   END n_35567

   PIN n_3607
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 64.15 0.51 64.25 ;
      END
   END n_3607

   PIN n_3623
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 12.75 0.51 12.85 ;
      END
   END n_3623

   PIN n_3863
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 10.55 0.51 10.65 ;
      END
   END n_3863

   PIN n_3903
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 6.45 0 6.55 0.51 ;
      END
   END n_3903

   PIN n_3909
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.65 0 8.75 0.51 ;
      END
   END n_3909

   PIN n_3935
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 10.35 0.51 10.45 ;
      END
   END n_3935

   PIN n_4062
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 3.65 0 3.75 0.51 ;
      END
   END n_4062

   PIN n_4064
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 64.35 0.51 64.45 ;
      END
   END n_4064

   PIN n_4068
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 26.15 0.51 26.25 ;
      END
   END n_4068

   PIN n_4079
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 10.15 0.51 10.25 ;
      END
   END n_4079

   PIN n_4088
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 12.85 0 12.95 0.51 ;
      END
   END n_4088

   PIN n_4104
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 20.75 0.51 20.85 ;
      END
   END n_4104

   PIN n_4105
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 28.85 0 28.95 0.51 ;
      END
   END n_4105

   PIN n_4118
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.15 0.51 33.25 ;
      END
   END n_4118

   PIN n_4122
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.05 0 31.15 0.51 ;
      END
   END n_4122

   PIN n_4131
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.25 0 19.35 0.51 ;
      END
   END n_4131

   PIN n_4201
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 64.55 0.51 64.65 ;
      END
   END n_4201

   PIN n_4204
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 30.85 0 30.95 0.51 ;
      END
   END n_4204

   PIN n_4294
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.45 0 3.55 0.51 ;
      END
   END n_4294

   PIN n_4490
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 7.45 0 7.55 0.51 ;
      END
   END n_4490

   PIN n_4494
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.25 0 8.35 0.51 ;
      END
   END n_4494

   PIN n_4561
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 1.25 0 1.35 0.51 ;
      END
   END n_4561

   PIN n_4708
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 34.45 0 34.55 0.51 ;
      END
   END n_4708

   PIN n_4799
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 11.55 0.51 11.65 ;
      END
   END n_4799

   PIN n_4811
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 5.25 0 5.35 0.51 ;
      END
   END n_4811

   PIN n_4882
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.95 0.51 22.05 ;
      END
   END n_4882

   PIN n_4923
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 9.05 0 9.15 0.51 ;
      END
   END n_4923

   PIN n_4958
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 25.65 0 25.75 0.51 ;
      END
   END n_4958

   PIN n_4961
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 50.15 0.51 50.25 ;
      END
   END n_4961

   PIN n_5049
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 50.35 0.51 50.45 ;
      END
   END n_5049

   PIN n_5069
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.25 0 33.35 0.51 ;
      END
   END n_5069

   PIN n_5268
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.45 0 23.55 0.51 ;
      END
   END n_5268

   PIN n_5314
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.25 0 31.35 0.51 ;
      END
   END n_5314

   PIN n_5323
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 41.45 0 41.55 0.51 ;
      END
   END n_5323

   PIN n_5363
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 24.45 0 24.55 0.51 ;
      END
   END n_5363

   PIN n_5372
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.55 0.51 75.65 ;
      END
   END n_5372

   PIN n_5437
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37.65 0 37.75 0.51 ;
      END
   END n_5437

   PIN n_5482
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.05 0 42.15 0.51 ;
      END
   END n_5482

   PIN n_5571
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.05 0 47.15 0.51 ;
      END
   END n_5571

   PIN n_5574
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 76.15 0.51 76.25 ;
      END
   END n_5574

   PIN n_5581
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 37.95 0.51 38.05 ;
      END
   END n_5581

   PIN n_5643
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.85 0 38.95 0.51 ;
      END
   END n_5643

   PIN n_59574
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 32.15 0.51 32.25 ;
      END
   END n_59574

   PIN n_6096
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.45 0 59.55 0.51 ;
      END
   END n_6096

   PIN n_61534
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 14.15 0.51 14.25 ;
      END
   END n_61534

   PIN n_61611
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 2.45 0 2.55 0.51 ;
      END
   END n_61611

   PIN n_6257
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 39.25 0 39.35 0.51 ;
      END
   END n_6257

   PIN n_63161
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.95 0.51 28.05 ;
      END
   END n_63161

   PIN n_63230
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 116.05 295.49 116.15 296 ;
      END
   END n_63230

   PIN n_63234
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.15 0.51 31.25 ;
      END
   END n_63234

   PIN n_63421
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 34.95 0.51 35.05 ;
      END
   END n_63421

   PIN n_63508
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 11.05 0 11.15 0.51 ;
      END
   END n_63508

   PIN n_63603
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.25 0 67.35 0.51 ;
      END
   END n_63603

   PIN n_63622
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 184.35 0.51 184.45 ;
      END
   END n_63622

   PIN n_63690
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 102.15 0.51 102.25 ;
      END
   END n_63690

   PIN n_63695
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.35 0.51 88.45 ;
      END
   END n_63695

   PIN n_63776
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 183.75 0.51 183.85 ;
      END
   END n_63776

   PIN n_63794
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 65.45 0 65.55 0.51 ;
      END
   END n_63794

   PIN n_63840
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 73.65 0 73.75 0.51 ;
      END
   END n_63840

   PIN n_63851
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.45 0 71.55 0.51 ;
      END
   END n_63851

   PIN n_63858
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.2 0 72.4 0.255 ;
      END
   END n_63858

   PIN n_63883
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.85 0 73.95 0.51 ;
      END
   END n_63883

   PIN n_63885
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 75.25 0 75.35 0.51 ;
      END
   END n_63885

   PIN n_63886
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.85 0 72.95 0.51 ;
      END
   END n_63886

   PIN n_63972
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 65.25 0 65.35 0.51 ;
      END
   END n_63972

   PIN n_64022
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.65 0 70.75 0.51 ;
      END
   END n_64022

   PIN n_64028
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 148.15 0.51 148.25 ;
      END
   END n_64028

   PIN n_64034
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.25 0 16.35 0.51 ;
      END
   END n_64034

   PIN n_64049
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.25 0 68.35 0.51 ;
      END
   END n_64049

   PIN n_64091
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 88.15 0.51 88.25 ;
      END
   END n_64091

   PIN n_64119
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 102.5 0.255 102.7 ;
      END
   END n_64119

   PIN n_64138
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.65 0 64.75 0.51 ;
      END
   END n_64138

   PIN n_64153
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 99.95 0.51 100.05 ;
      END
   END n_64153

   PIN n_64188
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 184.15 0.51 184.25 ;
      END
   END n_64188

   PIN n_64189
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 183.95 0.51 184.05 ;
      END
   END n_64189

   PIN n_64248
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.25 0 72.35 0.51 ;
      END
   END n_64248

   PIN n_64308
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 88.35 0.51 88.45 ;
      END
   END n_64308

   PIN n_64341
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 183.55 0.51 183.65 ;
      END
   END n_64341

   PIN n_64388
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 72.05 0 72.15 0.51 ;
      END
   END n_64388

   PIN n_64414
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 99.75 0.51 99.85 ;
      END
   END n_64414

   PIN n_64439
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 75.05 0 75.15 0.51 ;
      END
   END n_64439

   PIN n_64590
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.45 0 67.55 0.51 ;
      END
   END n_64590

   PIN n_64618
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.05 0 78.15 0.51 ;
      END
   END n_64618

   PIN n_64713
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.85 0 77.95 0.51 ;
      END
   END n_64713

   PIN n_64732
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.45 0 70.55 0.51 ;
      END
   END n_64732

   PIN n_64733
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.65 0 77.75 0.51 ;
      END
   END n_64733

   PIN n_64736
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.85 0 67.95 0.51 ;
      END
   END n_64736

   PIN n_64749
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.85 0 71.95 0.51 ;
      END
   END n_64749

   PIN n_64824
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 65.65 0 65.75 0.51 ;
      END
   END n_64824

   PIN n_64842
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.05 0 77.15 0.51 ;
      END
   END n_64842

   PIN n_64909
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 65.25 0 65.35 0.51 ;
      END
   END n_64909

   PIN n_64922
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 62.85 0 62.95 0.51 ;
      END
   END n_64922

   PIN n_64923
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 65.05 0 65.15 0.51 ;
      END
   END n_64923

   PIN n_64962
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 195.55 0.51 195.65 ;
      END
   END n_64962

   PIN n_65028
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 93.25 0 93.35 0.51 ;
      END
   END n_65028

   PIN n_6503
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 192.65 0 192.75 0.51 ;
      END
   END n_6503

   PIN n_65155
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.05 0 64.15 0.51 ;
      END
   END n_65155

   PIN n_65446
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.85 0 20.95 0.51 ;
      END
   END n_65446

   PIN n_65451
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 21.25 0 21.35 0.51 ;
      END
   END n_65451

   PIN n_65473
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.35 0.51 124.45 ;
      END
   END n_65473

   PIN n_65475
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 87.05 0 87.15 0.51 ;
      END
   END n_65475

   PIN n_65507
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.55 0.51 41.65 ;
      END
   END n_65507

   PIN n_65527
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.7 0.255 35.9 ;
      END
   END n_65527

   PIN n_65552
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 31.95 0.51 32.05 ;
      END
   END n_65552

   PIN n_65560
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.25 0 38.35 0.51 ;
      END
   END n_65560

   PIN n_65578
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.45 0 47.55 0.51 ;
      END
   END n_65578

   PIN n_65583
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 42.35 0.51 42.45 ;
      END
   END n_65583

   PIN n_65610
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.55 0.51 38.65 ;
      END
   END n_65610

   PIN n_65621
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 43.35 0.51 43.45 ;
      END
   END n_65621

   PIN n_65671
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 85.65 0 85.75 0.51 ;
      END
   END n_65671

   PIN n_65702
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.65 0 47.75 0.51 ;
      END
   END n_65702

   PIN n_65747
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.85 0 47.95 0.51 ;
      END
   END n_65747

   PIN n_65752
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 82.45 0 82.55 0.51 ;
      END
   END n_65752

   PIN n_65753
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 13.95 0.51 14.05 ;
      END
   END n_65753

   PIN n_65810
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.15 0.51 39.25 ;
      END
   END n_65810

   PIN n_65890
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.55 0.51 50.65 ;
      END
   END n_65890

   PIN n_65897
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.55 0.51 37.65 ;
      END
   END n_65897

   PIN n_65923
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 81.45 0 81.55 0.51 ;
      END
   END n_65923

   PIN n_65941
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.35 0.51 32.45 ;
      END
   END n_65941

   PIN n_65953
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.75 0.51 38.85 ;
      END
   END n_65953

   PIN n_65962
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 82.85 0 82.95 0.51 ;
      END
   END n_65962

   PIN n_65965
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 83.25 0 83.35 0.51 ;
      END
   END n_65965

   PIN n_65979
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.75 0.51 50.85 ;
      END
   END n_65979

   PIN n_66001
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 46.65 0 46.75 0.51 ;
      END
   END n_66001

   PIN n_66004
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44.45 0 44.55 0.51 ;
      END
   END n_66004

   PIN n_66070
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 85.85 0 85.95 0.51 ;
      END
   END n_66070

   PIN n_66106
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.15 0.51 38.25 ;
      END
   END n_66106

   PIN n_66122
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 50.45 0 50.55 0.51 ;
      END
   END n_66122

   PIN n_66130
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.55 0.51 51.65 ;
      END
   END n_66130

   PIN n_66184
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.85 0 80.95 0.51 ;
      END
   END n_66184

   PIN n_66209
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 81.25 0 81.35 0.51 ;
      END
   END n_66209

   PIN n_66223
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.85 0 81.95 0.51 ;
      END
   END n_66223

   PIN n_66292
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 84.65 0 84.75 0.51 ;
      END
   END n_66292

   PIN n_66319
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.05 295.49 128.15 296 ;
      END
   END n_66319

   PIN n_66357
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 45.05 0 45.15 0.51 ;
      END
   END n_66357

   PIN n_66374
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 79.6 0 79.8 0.255 ;
      END
   END n_66374

   PIN n_66380
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 12.55 0.51 12.65 ;
      END
   END n_66380

   PIN n_66389
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.05 0 80.15 0.51 ;
      END
   END n_66389

   PIN n_66417
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 50.75 0.51 50.85 ;
      END
   END n_66417

   PIN n_66438
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 12.35 0.51 12.45 ;
      END
   END n_66438

   PIN n_66469
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.05 0 81.15 0.51 ;
      END
   END n_66469

   PIN n_66475
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 42.45 0 42.55 0.51 ;
      END
   END n_66475

   PIN n_66487
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.35 0.51 35.45 ;
      END
   END n_66487

   PIN n_66506
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.05 0 91.15 0.51 ;
      END
   END n_66506

   PIN n_66569
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 40.65 0 40.75 0.51 ;
      END
   END n_66569

   PIN n_66584
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.65 0 43.75 0.51 ;
      END
   END n_66584

   PIN n_66589
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 42.05 0 42.15 0.51 ;
      END
   END n_66589

   PIN n_66623
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.35 0.51 37.45 ;
      END
   END n_66623

   PIN n_66630
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.15 0.51 37.25 ;
      END
   END n_66630

   PIN n_66656
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 99.55 0.51 99.65 ;
      END
   END n_66656

   PIN n_66678
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 45.45 0 45.55 0.51 ;
      END
   END n_66678

   PIN n_66807
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 0.85 0 0.95 0.51 ;
      END
   END n_66807

   PIN n_66822
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.75 0.51 111.85 ;
      END
   END n_66822

   PIN n_66873
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.95 0.51 37.05 ;
      END
   END n_66873

   PIN n_67053
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 32.75 0.51 32.85 ;
      END
   END n_67053

   PIN n_67065
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.85 295.49 127.95 296 ;
      END
   END n_67065

   PIN n_67119
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.75 0.51 36.85 ;
      END
   END n_67119

   PIN n_67131
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.45 295.49 56.55 296 ;
      END
   END n_67131

   PIN n_67150
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.15 0.51 124.25 ;
      END
   END n_67150

   PIN n_67203
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 10.55 0.51 10.65 ;
      END
   END n_67203

   PIN n_67231
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.95 0.51 124.05 ;
      END
   END n_67231

   PIN n_67232
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 123.75 0.51 123.85 ;
      END
   END n_67232

   PIN n_67245
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 132.05 295.49 132.15 296 ;
      END
   END n_67245

   PIN n_67246
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.45 295.49 127.55 296 ;
      END
   END n_67246

   PIN n_67247
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.05 295.49 116.15 296 ;
      END
   END n_67247

   PIN n_67326
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.05 295.49 56.15 296 ;
      END
   END n_67326

   PIN n_67480
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 58.05 0 58.15 0.51 ;
      END
   END n_67480

   PIN n_67630
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 54.2 0 54.4 0.255 ;
      END
   END n_67630

   PIN n_67644
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 54.85 0 54.95 0.51 ;
      END
   END n_67644

   PIN n_67654
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.65 0 48.75 0.51 ;
      END
   END n_67654

   PIN n_67771
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 58.25 0 58.35 0.51 ;
      END
   END n_67771

   PIN n_67793
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.05 0 56.15 0.51 ;
      END
   END n_67793

   PIN n_67946
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.25 0 52.35 0.51 ;
      END
   END n_67946

   PIN n_67996
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.85 0 126.95 0.51 ;
      END
   END n_67996

   PIN n_68009
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 53.85 0 53.95 0.51 ;
      END
   END n_68009

   PIN n_68020
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.15 0.51 88.25 ;
      END
   END n_68020

   PIN n_68045
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 57.45 0 57.55 0.51 ;
      END
   END n_68045

   PIN n_68057
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.95 0.51 88.05 ;
      END
   END n_68057

   PIN n_68205
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.45 0 48.55 0.51 ;
      END
   END n_68205

   PIN n_68264
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 90.85 0 90.95 0.51 ;
      END
   END n_68264

   PIN n_68269
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.05 0 52.15 0.51 ;
      END
   END n_68269

   PIN n_68283
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 54.25 0 54.35 0.51 ;
      END
   END n_68283

   PIN n_68286
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.85 0 48.95 0.51 ;
      END
   END n_68286

   PIN n_68349
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 78.45 0 78.55 0.51 ;
      END
   END n_68349

   PIN n_68352
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.25 0 56.35 0.51 ;
      END
   END n_68352

   PIN n_68366
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 54.65 0 54.75 0.51 ;
      END
   END n_68366

   PIN n_68377
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.85 0 59.95 0.51 ;
      END
   END n_68377

   PIN n_68515
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 47.25 0 47.35 0.51 ;
      END
   END n_68515

   PIN n_68805
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 53.65 0 53.75 0.51 ;
      END
   END n_68805

   PIN n_69023
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.95 0.51 76.05 ;
      END
   END n_69023

   PIN n_69052
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.75 0.51 75.85 ;
      END
   END n_69052

   PIN n_69101
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 87.75 0.51 87.85 ;
      END
   END n_69101

   PIN n_69155
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 49.75 0.51 49.85 ;
      END
   END n_69155

   PIN n_69285
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 38.55 0.51 38.65 ;
      END
   END n_69285

   PIN n_6944
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 92.25 0 92.35 0.51 ;
      END
   END n_6944

   PIN n_69515
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.25 0 55.35 0.51 ;
      END
   END n_69515

   PIN n_69551
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.35 0.51 51.45 ;
      END
   END n_69551

   PIN n_69624
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 66.05 0 66.15 0.51 ;
      END
   END n_69624

   PIN n_69650
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.65 0 36.75 0.51 ;
      END
   END n_69650

   PIN n_69668
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35.6 0 35.8 0.255 ;
      END
   END n_69668

   PIN n_69677
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.65 0 306.75 0.51 ;
      END
   END n_69677

   PIN n_69697
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 37.05 0 37.15 0.51 ;
      END
   END n_69697

   PIN n_69698
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.45 0 69.55 0.51 ;
      END
   END n_69698

   PIN n_69751
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 92.45 0 92.55 0.51 ;
      END
   END n_69751

   PIN n_69798
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 331.85 0 331.95 0.51 ;
      END
   END n_69798

   PIN n_69817
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.25 0 57.35 0.51 ;
      END
   END n_69817

   PIN n_69828
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 69.25 0 69.35 0.51 ;
      END
   END n_69828

   PIN n_69839
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 66.25 0 66.35 0.51 ;
      END
   END n_69839

   PIN n_70031
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.45 0 306.55 0.51 ;
      END
   END n_70031

   PIN n_70168
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 343.85 0 343.95 0.51 ;
      END
   END n_70168

   PIN n_70237
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 35.25 0 35.35 0.51 ;
      END
   END n_70237

   PIN n_70400
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 331.25 0 331.35 0.51 ;
      END
   END n_70400

   PIN n_70401
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 332.25 0 332.35 0.51 ;
      END
   END n_70401

   PIN n_70488
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 332.05 0 332.15 0.51 ;
      END
   END n_70488

   PIN n_70529
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 306.6 0 306.8 0.255 ;
      END
   END n_70529

   PIN n_70631
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.25 0 294.35 0.51 ;
      END
   END n_70631

   PIN n_70788
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.05 0 320.15 0.51 ;
      END
   END n_70788

   PIN n_7085
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 13.75 0.51 13.85 ;
      END
   END n_7085

   PIN n_70959
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 312.6 0 312.8 0.255 ;
      END
   END n_70959

   PIN n_70968
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.85 0 319.95 0.51 ;
      END
   END n_70968

   PIN n_70996
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 333.25 0 333.35 0.51 ;
      END
   END n_70996

   PIN n_71009
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 307.25 0 307.35 0.51 ;
      END
   END n_71009

   PIN n_71083
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.85 0 319.95 0.51 ;
      END
   END n_71083

   PIN n_71095
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 307.05 0 307.15 0.51 ;
      END
   END n_71095

   PIN n_71105
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.65 0 319.75 0.51 ;
      END
   END n_71105

   PIN n_71108
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 333.05 0 333.15 0.51 ;
      END
   END n_71108

   PIN n_71151
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.65 0 319.75 0.51 ;
      END
   END n_71151

   PIN n_71192
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.45 0 319.55 0.51 ;
      END
   END n_71192

   PIN n_7212
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 153.05 0 153.15 0.51 ;
      END
   END n_7212

   PIN n_753
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 38.35 0.51 38.45 ;
      END
   END n_753

   PIN n_75355
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.05 0 33.15 0.51 ;
      END
   END n_75355

   PIN n_75387
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 76.6 0 76.8 0.255 ;
      END
   END n_75387

   PIN n_75701
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 41.65 0 41.75 0.51 ;
      END
   END n_75701

   PIN n_75702
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 41.85 0 41.95 0.51 ;
      END
   END n_75702

   PIN n_75837
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.05 0 55.15 0.51 ;
      END
   END n_75837

   PIN n_75950
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 34.2 0 34.4 0.255 ;
      END
   END n_75950

   PIN n_75954
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 38.15 0.51 38.25 ;
      END
   END n_75954

   PIN n_76207
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 53.35 0.51 53.45 ;
      END
   END n_76207

   PIN n_76269
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 77.25 0 77.35 0.51 ;
      END
   END n_76269

   PIN n_76439
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 27.45 0 27.55 0.51 ;
      END
   END n_76439

   PIN n_76451
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 34.85 0 34.95 0.51 ;
      END
   END n_76451

   PIN n_76463
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 14.05 0 14.15 0.51 ;
      END
   END n_76463

   PIN n_76471
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 33.05 0 33.15 0.51 ;
      END
   END n_76471

   PIN n_76474
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 50.55 0.51 50.65 ;
      END
   END n_76474

   PIN n_76570
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.85 0 32.95 0.51 ;
      END
   END n_76570

   PIN n_76637
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.45 0 31.55 0.51 ;
      END
   END n_76637

   PIN n_76642
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 53.55 0.51 53.65 ;
      END
   END n_76642

   PIN n_76809
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 34.65 0 34.75 0.51 ;
      END
   END n_76809

   PIN n_76821
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 65.15 0.51 65.25 ;
      END
   END n_76821

   PIN n_77030
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 53.75 0.51 53.85 ;
      END
   END n_77030

   PIN n_77046
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 27.65 0 27.75 0.51 ;
      END
   END n_77046

   PIN n_77228
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 64.75 0.51 64.85 ;
      END
   END n_77228

   PIN n_77801
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 64.95 0.51 65.05 ;
      END
   END n_77801

   PIN n_78115
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 43.25 0 43.35 0.51 ;
      END
   END n_78115

   PIN n_7851
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.05 0 18.15 0.51 ;
      END
   END n_7851

   PIN n_7898
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 2.65 0 2.75 0.51 ;
      END
   END n_7898

   PIN n_90978
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 377.65 0 377.75 0.51 ;
      END
   END n_90978

   PIN n_95123
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 253.85 0 253.95 0.51 ;
      END
   END n_95123

   PIN n_9943
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.05 0 29.15 0.51 ;
      END
   END n_9943

   PIN stage1_out_3187
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 259.85 0 259.95 0.51 ;
      END
   END stage1_out_3187

   PIN stage1_out_3201
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 152.45 0 152.55 0.51 ;
      END
   END stage1_out_3201

   PIN stage1_out_3213
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 59.05 0 59.15 0.51 ;
      END
   END stage1_out_3213

   PIN u0_IP_64__1299
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.85 295.49 67.95 296 ;
      END
   END u0_IP_64__1299

   PIN u0_L4_29_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.95 0.51 35.05 ;
      END
   END u0_L4_29_

   PIN u0_L5_30_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 75.15 0.51 75.25 ;
      END
   END u0_L5_30_

   PIN u0_L6_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 24.95 0.51 25.05 ;
      END
   END u0_L6_10_

   PIN u0_L6_21_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.85 0 91.95 0.51 ;
      END
   END u0_L6_21_

   PIN u0_L6_29_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.05 0 140.15 0.51 ;
      END
   END u0_L6_29_

   PIN u0_L7_20_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 295.85 0 295.95 0.51 ;
      END
   END u0_L7_20_

   PIN u0_L7_28_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 152.85 0 152.95 0.51 ;
      END
   END u0_L7_28_

   PIN u0_L8_20_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 296.05 0 296.15 0.51 ;
      END
   END u0_L8_20_

   PIN u0_R2_26_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 21.15 0.51 21.25 ;
      END
   END u0_R2_26_

   PIN u0_R3_13_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 37.35 0.51 37.45 ;
      END
   END u0_R3_13_

   PIN u0_R3_16_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.65 0 163.75 0.51 ;
      END
   END u0_R3_16_

   PIN u0_R3_17_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.45 0 22.55 0.51 ;
      END
   END u0_R3_17_

   PIN u0_R3_19_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 49.35 0.51 49.45 ;
      END
   END u0_R3_19_

   PIN u0_R4_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 10.35 0.51 10.45 ;
      END
   END u0_R4_10_

   PIN u0_R4_17_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 74.95 0.51 75.05 ;
      END
   END u0_R4_17_

   PIN u0_R4_20_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 65.35 0.51 65.45 ;
      END
   END u0_R4_20_

   PIN u0_R5_13_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.25 295.49 56.35 296 ;
      END
   END u0_R5_13_

   PIN u0_R5_27_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 41.85 0 41.95 0.51 ;
      END
   END u0_R5_27_

   PIN u0_R5_4_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.05 295.49 20.15 296 ;
      END
   END u0_R5_4_

   PIN u0_R6_14_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 119.05 0 119.15 0.51 ;
      END
   END u0_R6_14_

   PIN u0_R6_17_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 49.55 0.51 49.65 ;
      END
   END u0_R6_17_

   PIN u0_R6_18_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 276.45 0 276.55 0.51 ;
      END
   END u0_R6_18_

   PIN u0_R6_23_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 313.45 0 313.55 0.51 ;
      END
   END u0_R6_23_

   PIN u0_R6_25_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 159.95 0.51 160.05 ;
      END
   END u0_R6_25_

   PIN u0_R6_26_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 367.05 0 367.15 0.51 ;
      END
   END u0_R6_26_

   PIN u0_R6_28_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 48.25 0 48.35 0.51 ;
      END
   END u0_R6_28_

   PIN u0_R6_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.05 0 63.15 0.51 ;
      END
   END u0_R6_3_

   PIN u0_R6_8_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 321.05 0 321.15 0.51 ;
      END
   END u0_R6_8_

   PIN u0_R7_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 201.65 0 201.75 0.51 ;
      END
   END u0_R7_10_

   PIN u0_R7_16_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 130.45 0 130.55 0.51 ;
      END
   END u0_R7_16_

   PIN u0_R7_20_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.25 0 197.35 0.51 ;
      END
   END u0_R7_20_

   PIN u0_R7_25_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 167.65 0 167.75 0.51 ;
      END
   END u0_R7_25_

   PIN u0_R7_28_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 120.65 0 120.75 0.51 ;
      END
   END u0_R7_28_

   PIN u0_R7_2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 194.65 0 194.75 0.51 ;
      END
   END u0_R7_2_

   PIN u0_R7_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 127.65 0 127.75 0.51 ;
      END
   END u0_R7_6_

   PIN u0_R8_23_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 301.45 0 301.55 0.51 ;
      END
   END u0_R8_23_

   PIN u0_key_r_23_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 115.05 0 115.15 0.51 ;
      END
   END u0_key_r_23_

   PIN u0_key_r_44_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.65 0 18.75 0.51 ;
      END
   END u0_key_r_44_

   PIN u0_uk_K_r_251
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 18.85 0 18.95 0.51 ;
      END
   END u0_uk_K_r_251

   PIN u0_uk_K_r_263
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.35 0.51 25.45 ;
      END
   END u0_uk_K_r_263

   PIN u0_uk_K_r_273
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.85 0 22.95 0.51 ;
      END
   END u0_uk_K_r_273

   PIN u0_uk_K_r_332
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.75 0.51 33.85 ;
      END
   END u0_uk_K_r_332

   PIN u0_uk_K_r_335
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 4.45 0 4.55 0.51 ;
      END
   END u0_uk_K_r_335

   PIN u0_uk_K_r_343
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 4.85 0 4.95 0.51 ;
      END
   END u0_uk_K_r_343

   PIN u0_uk_K_r_344
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 2.05 0 2.15 0.51 ;
      END
   END u0_uk_K_r_344

   PIN u0_uk_K_r_356
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.65 0 7.75 0.51 ;
      END
   END u0_uk_K_r_356

   PIN u0_uk_K_r_357
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 75.55 0.51 75.65 ;
      END
   END u0_uk_K_r_357

   PIN u0_uk_K_r_359
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 62.55 0.51 62.65 ;
      END
   END u0_uk_K_r_359

   PIN u0_uk_K_r_365
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 1.85 0 1.95 0.51 ;
      END
   END u0_uk_K_r_365

   PIN u0_uk_K_r_378
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.45 0 7.55 0.51 ;
      END
   END u0_uk_K_r_378

   PIN u0_uk_K_r_381
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.25 0 17.35 0.51 ;
      END
   END u0_uk_K_r_381

   PIN u0_uk_K_r_401
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.15 0.51 22.25 ;
      END
   END u0_uk_K_r_401

   PIN u0_uk_K_r_413
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 33.35 0.51 33.45 ;
      END
   END u0_uk_K_r_413

   PIN u0_uk_K_r_437
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 4.25 0 4.35 0.51 ;
      END
   END u0_uk_K_r_437

   PIN u0_uk_K_r_449
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 13.65 0 13.75 0.51 ;
      END
   END u0_uk_K_r_449

   PIN u0_uk_K_r_530
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 33.65 0 33.75 0.51 ;
      END
   END u0_uk_K_r_530

   PIN u1_L10_13_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.45 0 40.55 0.51 ;
      END
   END u1_L10_13_

   PIN u1_L11_22_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 37.15 0.51 37.25 ;
      END
   END u1_L11_22_

   PIN u1_L11_reg_7__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 47.75 0.51 47.85 ;
      END
   END u1_L11_reg_7__Q

   PIN u1_L7_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 36.75 0.51 36.85 ;
      END
   END u1_L7_7_

   PIN u1_R10_12_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.35 0.51 41.45 ;
      END
   END u1_R10_12_

   PIN u1_R8_19_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 41.15 0.51 41.25 ;
      END
   END u1_R8_19_

   PIN u1_R8_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 55.65 295.49 55.75 296 ;
      END
   END u1_R8_7_

   PIN u2_R6_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 309.05 0 309.15 0.51 ;
      END
   END u2_R6_7_

   PIN u2_R7_15_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.25 0 232.35 0.51 ;
      END
   END u2_R7_15_

   OBS
      LAYER via4 ;
         RECT 0 0 549.2 296 ;
      LAYER via3 ;
         RECT 0 0 549.2 296 ;
      LAYER via2 ;
         RECT 0 0 549.2 296 ;
      LAYER via1 ;
         RECT 0 0 549.2 296 ;
      LAYER metal5 ;
         RECT 0 0 549.2 296 ;
      LAYER metal4 ;
         RECT 0 0 549.2 296 ;
      LAYER metal3 ;
         RECT 0 0 549.2 296 ;
      LAYER metal2 ;
         RECT 0 0 549.2 296 ;
      LAYER metal1 ;
         RECT 0 0 549.2 296 ;
   END
END h3

MACRO h2
   CLASS BLOCK ;
   FOREIGN h2 ;
   ORIGIN 0 0 ;
   SIZE 523 BY 192 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1114_n_21429
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.25 191.49 161.35 192 ;
      END
   END FE_OFN1114_n_21429

   PIN FE_OFN1152_n_14527
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.45 191.49 291.55 192 ;
      END
   END FE_OFN1152_n_14527

   PIN FE_OFN1308_n_14014
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 210.85 191.49 210.95 192 ;
      END
   END FE_OFN1308_n_14014

   PIN FE_OFN13_n_106596
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 201.25 0 201.35 0.51 ;
      END
   END FE_OFN13_n_106596

   PIN FE_OFN1911_n_80620
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.65 191.49 103.75 192 ;
      END
   END FE_OFN1911_n_80620

   PIN FE_OFN194_n_84781
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.25 191.49 103.35 192 ;
      END
   END FE_OFN194_n_84781

   PIN FE_OFN200_n_15151
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.05 191.49 164.15 192 ;
      END
   END FE_OFN200_n_15151

   PIN FE_OFN2035_n_14525
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 166.45 191.49 166.55 192 ;
      END
   END FE_OFN2035_n_14525

   PIN FE_OFN2064_g190297_u0_o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 492.05 191.49 492.15 192 ;
      END
   END FE_OFN2064_g190297_u0_o

   PIN FE_OFN2073_n_107830
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 488.85 0 488.95 0.51 ;
      END
   END FE_OFN2073_n_107830

   PIN FE_OFN2234_n_75724
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 101.45 191.49 101.55 192 ;
      END
   END FE_OFN2234_n_75724

   PIN FE_OFN2250_n_82961
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 259.65 191.49 259.75 192 ;
      END
   END FE_OFN2250_n_82961

   PIN FE_OFN22_n_104304
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 288.45 191.49 288.55 192 ;
      END
   END FE_OFN22_n_104304

   PIN FE_OFN245_n_79557
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.85 191.49 199.95 192 ;
      END
   END FE_OFN245_n_79557

   PIN FE_OFN2549_n_118022
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 462.05 191.49 462.15 192 ;
      END
   END FE_OFN2549_n_118022

   PIN FE_OFN2763_n_107068
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 479.65 191.49 479.75 192 ;
      END
   END FE_OFN2763_n_107068

   PIN FE_OFN3492_n_83012
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 235.65 191.49 235.75 192 ;
      END
   END FE_OFN3492_n_83012

   PIN FE_OFN3552_n_81000
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 185.45 191.49 185.55 192 ;
      END
   END FE_OFN3552_n_81000

   PIN FE_OFN3554_n_108480
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 185.15 523 185.25 ;
      END
   END FE_OFN3554_n_108480

   PIN FE_OFN4785_n_77924
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.45 191.49 27.55 192 ;
      END
   END FE_OFN4785_n_77924

   PIN FE_OFN818_n_103115
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 236.85 191.49 236.95 192 ;
      END
   END FE_OFN818_n_103115

   PIN FE_OFN867_n_14026
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.25 191.49 116.35 192 ;
      END
   END FE_OFN867_n_14026

   PIN desOut_16_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 404.65 0 404.75 0.51 ;
      END
   END desOut_16_

   PIN desOut_17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 452.65 0 452.75 0.51 ;
      END
   END desOut_17_

   PIN desOut_38_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.65 0 128.75 0.51 ;
      END
   END desOut_38_

   PIN g190280_u0_o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 500.65 0 500.75 0.51 ;
      END
   END g190280_u0_o

   PIN g190611_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 462.25 191.49 462.35 192 ;
      END
   END g190611_p

   PIN g190906_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 47.95 523 48.05 ;
      END
   END g190906_p

   PIN g190953_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 154.95 523 155.05 ;
      END
   END g190953_p

   PIN g191131_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 155.75 523 155.85 ;
      END
   END g191131_p

   PIN g191163_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 155.15 523 155.25 ;
      END
   END g191163_p

   PIN g191647_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 380.45 191.49 380.55 192 ;
      END
   END g191647_da

   PIN g191647_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 375.65 191.49 375.75 192 ;
      END
   END g191647_db

   PIN g191648_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.05 0 163.15 0.51 ;
      END
   END g191648_da

   PIN g191648_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 172.45 0 172.55 0.51 ;
      END
   END g191648_db

   PIN g192426_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 358.25 191.49 358.35 192 ;
      END
   END g192426_p

   PIN g192601_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 187.65 191.49 187.75 192 ;
      END
   END g192601_p

   PIN g192862_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 81.95 0.51 82.05 ;
      END
   END g192862_p

   PIN g192893_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.15 0.51 71.25 ;
      END
   END g192893_p

   PIN g193052_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.65 0 224.75 0.51 ;
      END
   END g193052_p

   PIN g195141_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 150.45 191.49 150.55 192 ;
      END
   END g195141_da

   PIN g195175_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.05 191.49 283.15 192 ;
      END
   END g195175_p

   PIN g218222_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.25 191.49 291.35 192 ;
      END
   END g218222_sb

   PIN g218659_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 173.05 191.49 173.15 192 ;
      END
   END g218659_da

   PIN g218659_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 181.25 191.49 181.35 192 ;
      END
   END g218659_db

   PIN g219318_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 308.05 191.49 308.15 192 ;
      END
   END g219318_p

   PIN g219362_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 89.05 191.49 89.15 192 ;
      END
   END g219362_p

   PIN g219365_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 301.85 191.49 301.95 192 ;
      END
   END g219365_p

   PIN g220459_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 91.65 191.49 91.75 192 ;
      END
   END g220459_da

   PIN g220459_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.05 191.49 91.15 192 ;
      END
   END g220459_db

   PIN g223661_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 124.65 191.49 124.75 192 ;
      END
   END g223661_p

   PIN g223834_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 109.25 191.49 109.35 192 ;
      END
   END g223834_sb

   PIN g288188_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 227.05 191.49 227.15 192 ;
      END
   END g288188_p

   PIN g288202_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 217.45 191.49 217.55 192 ;
      END
   END g288202_p

   PIN g288612_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 79.65 191.49 79.75 192 ;
      END
   END g288612_p

   PIN key_c_r_31__2158
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 220.05 191.49 220.15 192 ;
      END
   END key_c_r_31__2158

   PIN key_c_r_33__8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 260.05 191.49 260.15 192 ;
      END
   END key_c_r_33__8_

   PIN n_100862
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 344.25 191.49 344.35 192 ;
      END
   END n_100862

   PIN n_100928
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 364.85 0 364.95 0.51 ;
      END
   END n_100928

   PIN n_101021
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 427.85 191.49 427.95 192 ;
      END
   END n_101021

   PIN n_102321
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 416.85 191.49 416.95 192 ;
      END
   END n_102321

   PIN n_102578
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 409.45 191.49 409.55 192 ;
      END
   END n_102578

   PIN n_103024
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 488.85 191.49 488.95 192 ;
      END
   END n_103024

   PIN n_103133
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 259.65 191.49 259.75 192 ;
      END
   END n_103133

   PIN n_103323
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 280.2 191.745 280.4 192 ;
      END
   END n_103323

   PIN n_103421
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.65 191.49 260.75 192 ;
      END
   END n_103421

   PIN n_103511
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.85 191.49 291.95 192 ;
      END
   END n_103511

   PIN n_103611
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 283.45 191.49 283.55 192 ;
      END
   END n_103611

   PIN n_103663
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 276.65 191.49 276.75 192 ;
      END
   END n_103663

   PIN n_103665
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 287.85 191.49 287.95 192 ;
      END
   END n_103665

   PIN n_103666
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 275.45 191.49 275.55 192 ;
      END
   END n_103666

   PIN n_103777
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.45 191.49 245.55 192 ;
      END
   END n_103777

   PIN n_103800
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 283.65 191.49 283.75 192 ;
      END
   END n_103800

   PIN n_103935
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.45 191.49 283.55 192 ;
      END
   END n_103935

   PIN n_104032
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 268.25 191.49 268.35 192 ;
      END
   END n_104032

   PIN n_104077
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 247.25 191.49 247.35 192 ;
      END
   END n_104077

   PIN n_104097
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 277.25 191.49 277.35 192 ;
      END
   END n_104097

   PIN n_104144
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.85 191.49 271.95 192 ;
      END
   END n_104144

   PIN n_104146
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 244.25 191.49 244.35 192 ;
      END
   END n_104146

   PIN n_104171
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 259.85 191.49 259.95 192 ;
      END
   END n_104171

   PIN n_104175
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 260.25 191.49 260.35 192 ;
      END
   END n_104175

   PIN n_104263
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 261.25 191.49 261.35 192 ;
      END
   END n_104263

   PIN n_104285
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 253.45 191.49 253.55 192 ;
      END
   END n_104285

   PIN n_104385
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.85 191.49 260.95 192 ;
      END
   END n_104385

   PIN n_104389
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 275.65 191.49 275.75 192 ;
      END
   END n_104389

   PIN n_104484
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 311.05 191.49 311.15 192 ;
      END
   END n_104484

   PIN n_104500
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.45 191.49 244.55 192 ;
      END
   END n_104500

   PIN n_104533
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 265.65 191.49 265.75 192 ;
      END
   END n_104533

   PIN n_104591
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.25 191.49 244.35 192 ;
      END
   END n_104591

   PIN n_104636
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 267.05 191.49 267.15 192 ;
      END
   END n_104636

   PIN n_104655
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 235.85 191.49 235.95 192 ;
      END
   END n_104655

   PIN n_104669
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.25 191.49 232.35 192 ;
      END
   END n_104669

   PIN n_105032
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 242.05 0 242.15 0.51 ;
      END
   END n_105032

   PIN n_105114
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 225 0 225.2 0.255 ;
      END
   END n_105114

   PIN n_105153
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 165.05 191.49 165.15 192 ;
      END
   END n_105153

   PIN n_105173
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 213.25 0 213.35 0.51 ;
      END
   END n_105173

   PIN n_105210
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 81.35 0.51 81.45 ;
      END
   END n_105210

   PIN n_105221
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.15 0.51 83.25 ;
      END
   END n_105221

   PIN n_105285
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.95 0.51 69.05 ;
      END
   END n_105285

   PIN n_105324
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 393.05 191.49 393.15 192 ;
      END
   END n_105324

   PIN n_105338
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 82.15 0.51 82.25 ;
      END
   END n_105338

   PIN n_105358
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.15 0.51 111.25 ;
      END
   END n_105358

   PIN n_105422
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.05 0 224.15 0.51 ;
      END
   END n_105422

   PIN n_105473
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 358.45 191.49 358.55 192 ;
      END
   END n_105473

   PIN n_105532
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.15 0.51 95.25 ;
      END
   END n_105532

   PIN n_105558
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.25 0 248.35 0.51 ;
      END
   END n_105558

   PIN n_105559
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 200.25 0 200.35 0.51 ;
      END
   END n_105559

   PIN n_105594
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.85 0 248.95 0.51 ;
      END
   END n_105594

   PIN n_105646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 200.05 0 200.15 0.51 ;
      END
   END n_105646

   PIN n_105647
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 215.05 0 215.15 0.51 ;
      END
   END n_105647

   PIN n_105690
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.65 0 164.75 0.51 ;
      END
   END n_105690

   PIN n_105698
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 370.05 191.49 370.15 192 ;
      END
   END n_105698

   PIN n_105744
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.25 0 212.35 0.51 ;
      END
   END n_105744

   PIN n_105750
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.05 0 188.15 0.51 ;
      END
   END n_105750

   PIN n_105751
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.65 0 248.75 0.51 ;
      END
   END n_105751

   PIN n_105789
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.55 0.51 52.65 ;
      END
   END n_105789

   PIN n_105899
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 59.95 0.51 60.05 ;
      END
   END n_105899

   PIN n_105911
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.25 0 188.35 0.51 ;
      END
   END n_105911

   PIN n_105913
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.65 0 176.75 0.51 ;
      END
   END n_105913

   PIN n_105936
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 181.25 0 181.35 0.51 ;
      END
   END n_105936

   PIN n_105940
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 242.2 0 242.4 0.255 ;
      END
   END n_105940

   PIN n_105951
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 61.15 0.51 61.25 ;
      END
   END n_105951

   PIN n_105999
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 369.85 191.49 369.95 192 ;
      END
   END n_105999

   PIN n_106024
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 353.85 191.49 353.95 192 ;
      END
   END n_106024

   PIN n_106031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.45 0 152.55 0.51 ;
      END
   END n_106031

   PIN n_106032
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 200.65 0 200.75 0.51 ;
      END
   END n_106032

   PIN n_106044
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 387.85 191.49 387.95 192 ;
      END
   END n_106044

   PIN n_106048
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.65 0 308.75 0.51 ;
      END
   END n_106048

   PIN n_106077
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 60.15 0.51 60.25 ;
      END
   END n_106077

   PIN n_106100
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.35 0.51 71.45 ;
      END
   END n_106100

   PIN n_106152
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 61.75 0.51 61.85 ;
      END
   END n_106152

   PIN n_106178
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.35 0.51 68.45 ;
      END
   END n_106178

   PIN n_106206
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 365.25 191.49 365.35 192 ;
      END
   END n_106206

   PIN n_106225
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 187.65 0 187.75 0.51 ;
      END
   END n_106225

   PIN n_106257
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 61.35 0.51 61.45 ;
      END
   END n_106257

   PIN n_106305
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 375.85 191.49 375.95 192 ;
      END
   END n_106305

   PIN n_106309
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 376.25 191.49 376.35 192 ;
      END
   END n_106309

   PIN n_106315
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 191.85 0 191.95 0.51 ;
      END
   END n_106315

   PIN n_106345
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 380.25 191.49 380.35 192 ;
      END
   END n_106345

   PIN n_106356
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.85 0 197.95 0.51 ;
      END
   END n_106356

   PIN n_106374
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.95 0.51 81.05 ;
      END
   END n_106374

   PIN n_106382
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 516.85 191.49 516.95 192 ;
      END
   END n_106382

   PIN n_106401
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 384.85 191.49 384.95 192 ;
      END
   END n_106401

   PIN n_106404
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.55 0.51 95.65 ;
      END
   END n_106404

   PIN n_106446
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.85 0 164.95 0.51 ;
      END
   END n_106446

   PIN n_106447
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.65 0 152.75 0.51 ;
      END
   END n_106447

   PIN n_106458
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 47.15 0.51 47.25 ;
      END
   END n_106458

   PIN n_106496
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 380.05 191.49 380.15 192 ;
      END
   END n_106496

   PIN n_106527
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.55 0.51 68.65 ;
      END
   END n_106527

   PIN n_106534
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.95 0.51 52.05 ;
      END
   END n_106534

   PIN n_106558
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 118.65 0 118.75 0.51 ;
      END
   END n_106558

   PIN n_106576
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 61.55 0.51 61.65 ;
      END
   END n_106576

   PIN n_106582
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 66.95 0.51 67.05 ;
      END
   END n_106582

   PIN n_106653
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 379.85 191.49 379.95 192 ;
      END
   END n_106653

   PIN n_106665
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.05 0 164.15 0.51 ;
      END
   END n_106665

   PIN n_106667
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.75 0.51 52.85 ;
      END
   END n_106667

   PIN n_106671
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 200.05 191.49 200.15 192 ;
      END
   END n_106671

   PIN n_106682
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 383.45 191.49 383.55 192 ;
      END
   END n_106682

   PIN n_106715
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.85 0 123.95 0.51 ;
      END
   END n_106715

   PIN n_106742
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 392.85 191.49 392.95 192 ;
      END
   END n_106742

   PIN n_106753
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 223.45 191.49 223.55 192 ;
      END
   END n_106753

   PIN n_106769
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.65 191.49 132.75 192 ;
      END
   END n_106769

   PIN n_106772
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 187.85 191.49 187.95 192 ;
      END
   END n_106772

   PIN n_106806
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 452.25 191.49 452.35 192 ;
      END
   END n_106806

   PIN n_106814
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.65 0 151.75 0.51 ;
      END
   END n_106814

   PIN n_106816
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.85 0 141.95 0.51 ;
      END
   END n_106816

   PIN n_106875
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.45 191.49 163.55 192 ;
      END
   END n_106875

   PIN n_107039
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 501.05 191.49 501.15 192 ;
      END
   END n_107039

   PIN n_107087
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 511.25 0 511.35 0.51 ;
      END
   END n_107087

   PIN n_107115
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 167.95 523 168.05 ;
      END
   END n_107115

   PIN n_107137
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 513.05 191.49 513.15 192 ;
      END
   END n_107137

   PIN n_107138
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 465.05 191.49 465.15 192 ;
      END
   END n_107138

   PIN n_107156
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 512.65 191.49 512.75 192 ;
      END
   END n_107156

   PIN n_107223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 475.65 191.49 475.75 192 ;
      END
   END n_107223

   PIN n_107261
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 464.05 191.49 464.15 192 ;
      END
   END n_107261

   PIN n_107361
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 512.85 191.49 512.95 192 ;
      END
   END n_107361

   PIN n_107390
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 477.25 191.49 477.35 192 ;
      END
   END n_107390

   PIN n_107391
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 475.85 191.49 475.95 192 ;
      END
   END n_107391

   PIN n_107409
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 499.25 0 499.35 0.51 ;
      END
   END n_107409

   PIN n_107414
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 464.45 191.49 464.55 192 ;
      END
   END n_107414

   PIN n_107424
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 509.65 0 509.75 0.51 ;
      END
   END n_107424

   PIN n_107426
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 452.05 0 452.15 0.51 ;
      END
   END n_107426

   PIN n_107429
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 36.95 523 37.05 ;
      END
   END n_107429

   PIN n_107430
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 500.45 0 500.55 0.51 ;
      END
   END n_107430

   PIN n_107482
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 464.65 191.49 464.75 192 ;
      END
   END n_107482

   PIN n_107485
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 143.75 523 143.85 ;
      END
   END n_107485

   PIN n_107498
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 512.65 0 512.75 0.51 ;
      END
   END n_107498

   PIN n_107515
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 464.85 191.49 464.95 192 ;
      END
   END n_107515

   PIN n_107520
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 488.05 191.49 488.15 192 ;
      END
   END n_107520

   PIN n_107556
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 81.35 523 81.45 ;
      END
   END n_107556

   PIN n_107586
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 11.95 523 12.05 ;
      END
   END n_107586

   PIN n_107658
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 500.85 0 500.95 0.51 ;
      END
   END n_107658

   PIN n_107704
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 80.95 523 81.05 ;
      END
   END n_107704

   PIN n_107733
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 500.65 191.49 500.75 192 ;
      END
   END n_107733

   PIN n_107740
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 392.45 0 392.55 0.51 ;
      END
   END n_107740

   PIN n_107831
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 510.25 0 510.35 0.51 ;
      END
   END n_107831

   PIN n_107875
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 464.45 191.49 464.55 192 ;
      END
   END n_107875

   PIN n_107879
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 496.65 0 496.75 0.51 ;
      END
   END n_107879

   PIN n_107901
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 476.65 0 476.75 0.51 ;
      END
   END n_107901

   PIN n_107909
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 476.45 191.49 476.55 192 ;
      END
   END n_107909

   PIN n_107910
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 469.25 0 469.35 0.51 ;
      END
   END n_107910

   PIN n_107929
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 500.65 191.49 500.75 192 ;
      END
   END n_107929

   PIN n_107930
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 466.05 191.49 466.15 192 ;
      END
   END n_107930

   PIN n_107938
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 483.65 191.49 483.75 192 ;
      END
   END n_107938

   PIN n_107997
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 488.45 191.49 488.55 192 ;
      END
   END n_107997

   PIN n_107998
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 451.85 0 451.95 0.51 ;
      END
   END n_107998

   PIN n_108000
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 119.95 523 120.05 ;
      END
   END n_108000

   PIN n_108052
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 513.25 191.49 513.35 192 ;
      END
   END n_108052

   PIN n_108056
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 487.8 191.745 488 192 ;
      END
   END n_108056

   PIN n_108058
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 464.25 191.49 464.35 192 ;
      END
   END n_108058

   PIN n_108059
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 463.85 191.49 463.95 192 ;
      END
   END n_108059

   PIN n_108064
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 503.65 0 503.75 0.51 ;
      END
   END n_108064

   PIN n_108065
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 83.55 523 83.65 ;
      END
   END n_108065

   PIN n_108083
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 460.05 191.49 460.15 192 ;
      END
   END n_108083

   PIN n_108088
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 488.65 0 488.75 0.51 ;
      END
   END n_108088

   PIN n_108129
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 50.95 523 51.05 ;
      END
   END n_108129

   PIN n_108132
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 502.65 0 502.75 0.51 ;
      END
   END n_108132

   PIN n_108133
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 467.45 0 467.55 0.51 ;
      END
   END n_108133

   PIN n_108161
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 475.45 191.49 475.55 192 ;
      END
   END n_108161

   PIN n_108172
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 477.05 191.49 477.15 192 ;
      END
   END n_108172

   PIN n_108179
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 448.25 191.49 448.35 192 ;
      END
   END n_108179

   PIN n_108192
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 446.85 191.49 446.95 192 ;
      END
   END n_108192

   PIN n_108216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 72.15 523 72.25 ;
      END
   END n_108216

   PIN n_108224
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 500.85 191.49 500.95 192 ;
      END
   END n_108224

   PIN n_108227
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 83.95 523 84.05 ;
      END
   END n_108227

   PIN n_108234
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 476.85 191.49 476.95 192 ;
      END
   END n_108234

   PIN n_108235
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 476.65 191.49 476.75 192 ;
      END
   END n_108235

   PIN n_108244
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 125.15 523 125.25 ;
      END
   END n_108244

   PIN n_108274
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 513.45 191.49 513.55 192 ;
      END
   END n_108274

   PIN n_108297
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 184.95 523 185.05 ;
      END
   END n_108297

   PIN n_108300
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 476.85 191.49 476.95 192 ;
      END
   END n_108300

   PIN n_108311
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 476.05 191.49 476.15 192 ;
      END
   END n_108311

   PIN n_108318
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 477.45 191.49 477.55 192 ;
      END
   END n_108318

   PIN n_108320
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 477.45 191.49 477.55 192 ;
      END
   END n_108320

   PIN n_108329
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 477.05 191.49 477.15 192 ;
      END
   END n_108329

   PIN n_108337
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 185.35 523 185.45 ;
      END
   END n_108337

   PIN n_108392
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 155.35 523 155.45 ;
      END
   END n_108392

   PIN n_108450
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 477.65 191.49 477.75 192 ;
      END
   END n_108450

   PIN n_108486
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 475.05 191.49 475.15 192 ;
      END
   END n_108486

   PIN n_112858
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 249.25 191.49 249.35 192 ;
      END
   END n_112858

   PIN n_112987
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 462.65 0 462.75 0.51 ;
      END
   END n_112987

   PIN n_117115
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.85 191.49 255.95 192 ;
      END
   END n_117115

   PIN n_118365
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 288.25 191.49 288.35 192 ;
      END
   END n_118365

   PIN n_118376
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 277.45 191.49 277.55 192 ;
      END
   END n_118376

   PIN n_118637
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 380.25 191.49 380.35 192 ;
      END
   END n_118637

   PIN n_126056
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 337.45 191.49 337.55 192 ;
      END
   END n_126056

   PIN n_126215
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 36.95 0.51 37.05 ;
      END
   END n_126215

   PIN n_13159
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.05 191.49 140.15 192 ;
      END
   END n_13159

   PIN n_13183
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 117.65 191.49 117.75 192 ;
      END
   END n_13183

   PIN n_13379
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.65 191.49 91.75 192 ;
      END
   END n_13379

   PIN n_13383
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 145.25 191.49 145.35 192 ;
      END
   END n_13383

   PIN n_13413
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 224.05 191.49 224.15 192 ;
      END
   END n_13413

   PIN n_13426
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 103.25 191.49 103.35 192 ;
      END
   END n_13426

   PIN n_13478
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 89.45 191.49 89.55 192 ;
      END
   END n_13478

   PIN n_13607
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.05 191.49 112.15 192 ;
      END
   END n_13607

   PIN n_13698
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 117.05 191.49 117.15 192 ;
      END
   END n_13698

   PIN n_137144
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.95 0.51 24.05 ;
      END
   END n_137144

   PIN n_137150
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.15 0.51 37.25 ;
      END
   END n_137150

   PIN n_13862
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 147.85 191.49 147.95 192 ;
      END
   END n_13862

   PIN n_13873
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 221.85 191.49 221.95 192 ;
      END
   END n_13873

   PIN n_13932
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 208.05 191.49 208.15 192 ;
      END
   END n_13932

   PIN n_14044
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.65 191.49 211.75 192 ;
      END
   END n_14044

   PIN n_14147
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.85 191.49 197.95 192 ;
      END
   END n_14147

   PIN n_14374
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 157.05 191.49 157.15 192 ;
      END
   END n_14374

   PIN n_14380
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 150.65 191.49 150.75 192 ;
      END
   END n_14380

   PIN n_183945
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.45 191.49 104.55 192 ;
      END
   END n_183945

   PIN n_183950
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 66.95 523 67.05 ;
      END
   END n_183950

   PIN n_75398
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 123.25 191.49 123.35 192 ;
      END
   END n_75398

   PIN n_75503
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.65 191.49 106.75 192 ;
      END
   END n_75503

   PIN n_75797
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 79.85 191.49 79.95 192 ;
      END
   END n_75797

   PIN n_75845
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.65 191.49 80.75 192 ;
      END
   END n_75845

   PIN n_75864
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.25 191.49 283.35 192 ;
      END
   END n_75864

   PIN n_75994
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 118.85 191.49 118.95 192 ;
      END
   END n_75994

   PIN n_76007
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 501.85 191.49 501.95 192 ;
      END
   END n_76007

   PIN n_76135
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.05 191.49 67.15 192 ;
      END
   END n_76135

   PIN n_76204
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 117.45 191.49 117.55 192 ;
      END
   END n_76204

   PIN n_76218
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 200.25 191.49 200.35 192 ;
      END
   END n_76218

   PIN n_76344
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 403.85 191.49 403.95 192 ;
      END
   END n_76344

   PIN n_76528
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 67.85 191.49 67.95 192 ;
      END
   END n_76528

   PIN n_76756
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 45.85 191.49 45.95 192 ;
      END
   END n_76756

   PIN n_76912
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 42.05 191.49 42.15 192 ;
      END
   END n_76912

   PIN n_76917
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.45 191.49 78.55 192 ;
      END
   END n_76917

   PIN n_76933
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 63.05 191.49 63.15 192 ;
      END
   END n_76933

   PIN n_76936
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 19.45 191.49 19.55 192 ;
      END
   END n_76936

   PIN n_76947
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 68.05 191.49 68.15 192 ;
      END
   END n_76947

   PIN n_76948
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 84.85 191.49 84.95 192 ;
      END
   END n_76948

   PIN n_76988
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.65 191.49 56.75 192 ;
      END
   END n_76988

   PIN n_77102
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 45.45 191.49 45.55 192 ;
      END
   END n_77102

   PIN n_77104
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 2.85 191.49 2.95 192 ;
      END
   END n_77104

   PIN n_77105
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.65 191.49 32.75 192 ;
      END
   END n_77105

   PIN n_77161
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.05 191.49 32.15 192 ;
      END
   END n_77161

   PIN n_77283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.05 191.49 3.15 192 ;
      END
   END n_77283

   PIN n_77379
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 50.25 191.49 50.35 192 ;
      END
   END n_77379

   PIN n_77468
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 32.05 191.49 32.15 192 ;
      END
   END n_77468

   PIN n_77547
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 7.25 191.49 7.35 192 ;
      END
   END n_77547

   PIN n_77747
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.25 191.49 44.35 192 ;
      END
   END n_77747

   PIN n_77781
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.85 191.49 32.95 192 ;
      END
   END n_77781

   PIN n_77819
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.25 191.49 32.35 192 ;
      END
   END n_77819

   PIN n_78099
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 23.85 191.49 23.95 192 ;
      END
   END n_78099

   PIN n_78517
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.25 191.49 16.35 192 ;
      END
   END n_78517

   PIN n_78714
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 85.25 191.49 85.35 192 ;
      END
   END n_78714

   PIN n_78796
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 70.65 191.49 70.75 192 ;
      END
   END n_78796

   PIN n_78872
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 71.65 191.49 71.75 192 ;
      END
   END n_78872

   PIN n_78903
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.85 191.49 185.95 192 ;
      END
   END n_78903

   PIN n_78996
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 223.65 191.49 223.75 192 ;
      END
   END n_78996

   PIN n_79015
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 415.05 191.49 415.15 192 ;
      END
   END n_79015

   PIN n_79054
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 425.05 191.49 425.15 192 ;
      END
   END n_79054

   PIN n_79058
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 416.05 191.49 416.15 192 ;
      END
   END n_79058

   PIN n_79069
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 237.45 191.49 237.55 192 ;
      END
   END n_79069

   PIN n_79114
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 97.65 191.49 97.75 192 ;
      END
   END n_79114

   PIN n_79207
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 337 191.745 337.2 192 ;
      END
   END n_79207

   PIN n_79217
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 439.25 191.49 439.35 192 ;
      END
   END n_79217

   PIN n_79224
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 440.65 191.49 440.75 192 ;
      END
   END n_79224

   PIN n_79290
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 117.45 191.49 117.55 192 ;
      END
   END n_79290

   PIN n_79306
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 118.2 191.745 118.4 192 ;
      END
   END n_79306

   PIN n_79355
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 431.85 191.49 431.95 192 ;
      END
   END n_79355

   PIN n_79357
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 428.25 191.49 428.35 192 ;
      END
   END n_79357

   PIN n_79378
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 438.85 191.49 438.95 192 ;
      END
   END n_79378

   PIN n_79379
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 442.65 191.49 442.75 192 ;
      END
   END n_79379

   PIN n_79388
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 181.85 191.49 181.95 192 ;
      END
   END n_79388

   PIN n_79399
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 422.65 191.49 422.75 192 ;
      END
   END n_79399

   PIN n_79410
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.85 191.49 103.95 192 ;
      END
   END n_79410

   PIN n_79432
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 335.05 191.49 335.15 192 ;
      END
   END n_79432

   PIN n_79456
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 105.05 191.49 105.15 192 ;
      END
   END n_79456

   PIN n_79462
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 439.65 191.49 439.75 192 ;
      END
   END n_79462

   PIN n_79483
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 413.05 191.49 413.15 192 ;
      END
   END n_79483

   PIN n_79497
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 248.65 191.49 248.75 192 ;
      END
   END n_79497

   PIN n_79507
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.05 191.49 152.15 192 ;
      END
   END n_79507

   PIN n_79513
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 128.8 191.745 129 192 ;
      END
   END n_79513

   PIN n_79516
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 179.25 191.49 179.35 192 ;
      END
   END n_79516

   PIN n_79537
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.25 191.49 140.35 192 ;
      END
   END n_79537

   PIN n_79569
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 184.65 191.49 184.75 192 ;
      END
   END n_79569

   PIN n_79577
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 148.2 191.745 148.4 192 ;
      END
   END n_79577

   PIN n_79626
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 200.65 191.49 200.75 192 ;
      END
   END n_79626

   PIN n_79648
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 276.8 191.745 277 192 ;
      END
   END n_79648

   PIN n_79650
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 404.05 191.49 404.15 192 ;
      END
   END n_79650

   PIN n_79680
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 237.85 191.49 237.95 192 ;
      END
   END n_79680

   PIN n_79682
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 127.65 191.49 127.75 192 ;
      END
   END n_79682

   PIN n_79688
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 177.25 191.49 177.35 192 ;
      END
   END n_79688

   PIN n_79690
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 109.05 191.49 109.15 192 ;
      END
   END n_79690

   PIN n_79712
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 415.85 191.49 415.95 192 ;
      END
   END n_79712

   PIN n_79715
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.05 191.49 104.15 192 ;
      END
   END n_79715

   PIN n_79718
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 345.65 0 345.75 0.51 ;
      END
   END n_79718

   PIN n_79779
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 437.45 191.49 437.55 192 ;
      END
   END n_79779

   PIN n_79782
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 427.65 191.49 427.75 192 ;
      END
   END n_79782

   PIN n_79783
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 415.65 191.49 415.75 192 ;
      END
   END n_79783

   PIN n_79785
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 423.05 191.49 423.15 192 ;
      END
   END n_79785

   PIN n_79863
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 247.45 191.49 247.55 192 ;
      END
   END n_79863

   PIN n_79879
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.05 191.49 92.15 192 ;
      END
   END n_79879

   PIN n_79888
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 165.25 191.49 165.35 192 ;
      END
   END n_79888

   PIN n_79920
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 416.65 191.49 416.75 192 ;
      END
   END n_79920

   PIN n_79923
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 417.25 191.49 417.35 192 ;
      END
   END n_79923

   PIN n_79934
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 428.45 191.49 428.55 192 ;
      END
   END n_79934

   PIN n_79946
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 188.05 191.49 188.15 192 ;
      END
   END n_79946

   PIN n_79982
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.25 0 293.35 0.51 ;
      END
   END n_79982

   PIN n_79989
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 339.05 191.49 339.15 192 ;
      END
   END n_79989

   PIN n_80001
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 142.45 191.49 142.55 192 ;
      END
   END n_80001

   PIN n_80015
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285.45 191.49 285.55 192 ;
      END
   END n_80015

   PIN n_80058
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 436.85 191.49 436.95 192 ;
      END
   END n_80058

   PIN n_80061
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 446.25 191.49 446.35 192 ;
      END
   END n_80061

   PIN n_80062
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 417.05 191.49 417.15 192 ;
      END
   END n_80062

   PIN n_80214
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 427.85 191.49 427.95 192 ;
      END
   END n_80214

   PIN n_80220
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 283.25 191.49 283.35 192 ;
      END
   END n_80220

   PIN n_80221
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 247.65 191.49 247.75 192 ;
      END
   END n_80221

   PIN n_80223
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 296.45 0 296.55 0.51 ;
      END
   END n_80223

   PIN n_80226
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 427.45 191.49 427.55 192 ;
      END
   END n_80226

   PIN n_80246
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 428.05 191.49 428.15 192 ;
      END
   END n_80246

   PIN n_80251
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.45 191.49 140.55 192 ;
      END
   END n_80251

   PIN n_80267
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.85 191.49 104.95 192 ;
      END
   END n_80267

   PIN n_80270
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 408.05 191.49 408.15 192 ;
      END
   END n_80270

   PIN n_80310
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.25 191.49 104.35 192 ;
      END
   END n_80310

   PIN n_80338
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 428.65 191.49 428.75 192 ;
      END
   END n_80338

   PIN n_80339
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 439.85 191.49 439.95 192 ;
      END
   END n_80339

   PIN n_80391
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 127.85 191.49 127.95 192 ;
      END
   END n_80391

   PIN n_80400
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.85 191.49 104.95 192 ;
      END
   END n_80400

   PIN n_80415
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 404.05 191.49 404.15 192 ;
      END
   END n_80415

   PIN n_80418
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 440.05 191.49 440.15 192 ;
      END
   END n_80418

   PIN n_80430
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 451.25 191.49 451.35 192 ;
      END
   END n_80430

   PIN n_80431
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 440.25 191.49 440.35 192 ;
      END
   END n_80431

   PIN n_80488
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 103.65 191.49 103.75 192 ;
      END
   END n_80488

   PIN n_80498
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 422.05 191.49 422.15 192 ;
      END
   END n_80498

   PIN n_80510
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.45 0 260.55 0.51 ;
      END
   END n_80510

   PIN n_80531
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 136.25 191.49 136.35 192 ;
      END
   END n_80531

   PIN n_80539
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 423.65 191.49 423.75 192 ;
      END
   END n_80539

   PIN n_80547
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.85 191.49 139.95 192 ;
      END
   END n_80547

   PIN n_80556
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 308.25 191.49 308.35 192 ;
      END
   END n_80556

   PIN n_80583
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.45 191.49 113.55 192 ;
      END
   END n_80583

   PIN n_80588
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 336.65 191.49 336.75 192 ;
      END
   END n_80588

   PIN n_80590
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 248.85 191.49 248.95 192 ;
      END
   END n_80590

   PIN n_80591
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.45 191.49 279.55 192 ;
      END
   END n_80591

   PIN n_80614
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.65 0 260.75 0.51 ;
      END
   END n_80614

   PIN n_80628
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.25 0 255.35 0.51 ;
      END
   END n_80628

   PIN n_80639
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 407.85 191.49 407.95 192 ;
      END
   END n_80639

   PIN n_80697
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 252.25 191.49 252.35 192 ;
      END
   END n_80697

   PIN n_80699
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 328.45 191.49 328.55 192 ;
      END
   END n_80699

   PIN n_80702
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 103.45 191.49 103.55 192 ;
      END
   END n_80702

   PIN n_80790
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.45 191.49 100.55 192 ;
      END
   END n_80790

   PIN n_80811
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.05 191.49 105.15 192 ;
      END
   END n_80811

   PIN n_80846
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 179.85 191.49 179.95 192 ;
      END
   END n_80846

   PIN n_80849
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.25 191.49 321.35 192 ;
      END
   END n_80849

   PIN n_80852
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 211.45 191.49 211.55 192 ;
      END
   END n_80852

   PIN n_80863
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 201.25 191.49 201.35 192 ;
      END
   END n_80863

   PIN n_80893
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 176.65 191.49 176.75 192 ;
      END
   END n_80893

   PIN n_81063
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 35.15 0.51 35.25 ;
      END
   END n_81063

   PIN n_81066
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 310.25 191.49 310.35 192 ;
      END
   END n_81066

   PIN n_81087
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 452.45 191.49 452.55 192 ;
      END
   END n_81087

   PIN n_81098
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.65 191.49 163.75 192 ;
      END
   END n_81098

   PIN n_81123
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.15 0.51 52.25 ;
      END
   END n_81123

   PIN n_81247
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 50.95 0.51 51.05 ;
      END
   END n_81247

   PIN n_81358
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 21.95 0.51 22.05 ;
      END
   END n_81358

   PIN n_81557
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 36.95 0.51 37.05 ;
      END
   END n_81557

   PIN n_81575
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 332.65 191.49 332.75 192 ;
      END
   END n_81575

   PIN n_81588
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.05 191.49 244.15 192 ;
      END
   END n_81588

   PIN n_81589
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 243.85 191.49 243.95 192 ;
      END
   END n_81589

   PIN n_81643
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 261.25 191.49 261.35 192 ;
      END
   END n_81643

   PIN n_81647
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 310.65 191.49 310.75 192 ;
      END
   END n_81647

   PIN n_81691
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.15 0.51 39.25 ;
      END
   END n_81691

   PIN n_81748
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 101.85 191.49 101.95 192 ;
      END
   END n_81748

   PIN n_81769
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 228.65 191.49 228.75 192 ;
      END
   END n_81769

   PIN n_81897
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.35 0.51 38.45 ;
      END
   END n_81897

   PIN n_81902
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 333.85 191.49 333.95 192 ;
      END
   END n_81902

   PIN n_81922
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 82.75 0.51 82.85 ;
      END
   END n_81922

   PIN n_81929
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.45 0 56.55 0.51 ;
      END
   END n_81929

   PIN n_81945
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.15 0.51 24.25 ;
      END
   END n_81945

   PIN n_81985
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 297.85 191.49 297.95 192 ;
      END
   END n_81985

   PIN n_82008
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 331.05 191.49 331.15 192 ;
      END
   END n_82008

   PIN n_82020
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.95 0.51 53.05 ;
      END
   END n_82020

   PIN n_82088
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 47.95 0.51 48.05 ;
      END
   END n_82088

   PIN n_82097
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 323.85 191.49 323.95 192 ;
      END
   END n_82097

   PIN n_82121
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.75 0.51 24.85 ;
      END
   END n_82121

   PIN n_82123
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.05 191.49 80.15 192 ;
      END
   END n_82123

   PIN n_82211
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 297.65 191.49 297.75 192 ;
      END
   END n_82211

   PIN n_82213
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 269.05 191.49 269.15 192 ;
      END
   END n_82213

   PIN n_82220
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 284.65 191.49 284.75 192 ;
      END
   END n_82220

   PIN n_82255
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.95 0.51 23.05 ;
      END
   END n_82255

   PIN n_82257
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.95 0.51 35.05 ;
      END
   END n_82257

   PIN n_82288
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.35 0.51 7.45 ;
      END
   END n_82288

   PIN n_82318
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 271.65 191.49 271.75 192 ;
      END
   END n_82318

   PIN n_82322
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 283.85 191.49 283.95 192 ;
      END
   END n_82322

   PIN n_82361
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.15 0.51 51.25 ;
      END
   END n_82361

   PIN n_82385
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 46.95 0.51 47.05 ;
      END
   END n_82385

   PIN n_82411
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 242.05 191.49 242.15 192 ;
      END
   END n_82411

   PIN n_82502
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.65 191.49 272.75 192 ;
      END
   END n_82502

   PIN n_82519
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 82.35 0.51 82.45 ;
      END
   END n_82519

   PIN n_82533
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 111.35 0.51 111.45 ;
      END
   END n_82533

   PIN n_82546
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285.85 191.49 285.95 192 ;
      END
   END n_82546

   PIN n_82552
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 316.85 191.49 316.95 192 ;
      END
   END n_82552

   PIN n_82605
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.35 0.51 52.45 ;
      END
   END n_82605

   PIN n_82608
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.45 191.49 320.55 192 ;
      END
   END n_82608

   PIN n_82617
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.85 191.49 91.95 192 ;
      END
   END n_82617

   PIN n_82646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 81.55 0.51 81.65 ;
      END
   END n_82646

   PIN n_82651
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.65 191.49 63.75 192 ;
      END
   END n_82651

   PIN n_82652
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 63.45 191.49 63.55 192 ;
      END
   END n_82652

   PIN n_82657
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.75 0.51 95.85 ;
      END
   END n_82657

   PIN n_82727
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.25 191.49 177.35 192 ;
      END
   END n_82727

   PIN n_82772
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 359.05 0 359.15 0.51 ;
      END
   END n_82772

   PIN n_82856
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 187.85 191.49 187.95 192 ;
      END
   END n_82856

   PIN n_82929
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.65 191.49 20.75 192 ;
      END
   END n_82929

   PIN n_82932
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.25 191.49 212.35 192 ;
      END
   END n_82932

   PIN n_82973
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 456.65 191.49 456.75 192 ;
      END
   END n_82973

   PIN n_83218
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 451.85 191.49 451.95 192 ;
      END
   END n_83218

   PIN n_83282
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 224.45 191.49 224.55 192 ;
      END
   END n_83282

   PIN n_83405
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 477.25 191.49 477.35 192 ;
      END
   END n_83405

   PIN n_83632
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 440.85 191.49 440.95 192 ;
      END
   END n_83632

   PIN stage2_out_3251
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 64.45 191.49 64.55 192 ;
      END
   END stage2_out_3251

   PIN stage2_out_3285
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 223.85 191.49 223.95 192 ;
      END
   END stage2_out_3285

   PIN u1_L14_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 200.45 191.49 200.55 192 ;
      END
   END u1_L14_6_

   PIN u1_L14_reg_29__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 91.05 191.49 91.15 192 ;
      END
   END u1_L14_reg_29__Q

   PIN u2_IP_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 49.05 191.49 49.15 192 ;
      END
   END u2_IP_1_

   PIN u2_IP_64__1283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.85 191.49 79.95 192 ;
      END
   END u2_IP_64__1283

   PIN u2_IP_64__1287
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 97.05 191.49 97.15 192 ;
      END
   END u2_IP_64__1287

   PIN u2_IP_64__1290
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.25 191.49 128.35 192 ;
      END
   END u2_IP_64__1290

   PIN u2_L0_21_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 356.25 191.49 356.35 192 ;
      END
   END u2_L0_21_

   PIN u2_L0_22_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 36.85 191.49 36.95 192 ;
      END
   END u2_L0_22_

   PIN u2_L12_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 371.85 191.49 371.95 192 ;
      END
   END u2_L12_15_

   PIN u2_L12_21_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 349.25 191.49 349.35 192 ;
      END
   END u2_L12_21_

   PIN u2_L12_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 344.45 191.49 344.55 192 ;
      END
   END u2_L12_5_

   PIN u2_L13_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 48.15 0.51 48.25 ;
      END
   END u2_L13_23_

   PIN u2_L13_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.65 0 139.75 0.51 ;
      END
   END u2_L13_28_

   PIN u2_L1_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 96.65 191.49 96.75 192 ;
      END
   END u2_L1_14_

   PIN u2_L1_25_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 103.85 191.49 103.95 192 ;
      END
   END u2_L1_25_

   PIN u2_L2_reg_7__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 223.45 191.49 223.55 192 ;
      END
   END u2_L2_reg_7__Q

   PIN u2_R0_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 151.85 191.49 151.95 192 ;
      END
   END u2_R0_28_

   PIN u2_R0_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 74.05 191.49 74.15 192 ;
      END
   END u2_R0_8_

   PIN u2_R11_5_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 236.45 191.49 236.55 192 ;
      END
   END u2_R11_5_

   PIN u2_R12_31_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.25 191.49 140.35 192 ;
      END
   END u2_R12_31_

   PIN u2_R13_15_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 489.05 191.49 489.15 192 ;
      END
   END u2_R13_15_

   PIN u2_R13_27_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 368.25 191.49 368.35 192 ;
      END
   END u2_R13_27_

   PIN u2_R14_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 488.25 191.49 488.35 192 ;
      END
   END u2_R14_6_

   PIN u2_R1_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 195.45 191.49 195.55 192 ;
      END
   END u2_R1_12_

   PIN u2_R1_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 235.45 191.49 235.55 192 ;
      END
   END u2_R1_7_

   PIN u2_R2_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.45 191.49 127.55 192 ;
      END
   END u2_R2_14_

   PIN u2_R2_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.65 191.49 44.75 192 ;
      END
   END u2_R2_23_

   PIN u2_R2_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 236.05 191.49 236.15 192 ;
      END
   END u2_R2_28_

   PIN u2_R3_11_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.85 0 283.95 0.51 ;
      END
   END u2_R3_11_

   PIN u2_R3_18_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 389.65 0 389.75 0.51 ;
      END
   END u2_R3_18_

   PIN u2_desIn_r_reg_12__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.25 191.49 71.35 192 ;
      END
   END u2_desIn_r_reg_12__Q

   PIN u2_key_r_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.45 191.49 163.55 192 ;
      END
   END u2_key_r_14_

   PIN u2_key_r_30_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.25 191.49 163.35 192 ;
      END
   END u2_key_r_30_

   PIN u2_key_r_43_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 211.65 191.49 211.75 192 ;
      END
   END u2_key_r_43_

   PIN u2_uk_K_r_222
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.85 191.49 139.95 192 ;
      END
   END u2_uk_K_r_222

   PIN u2_uk_K_r_365
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.25 191.49 92.35 192 ;
      END
   END u2_uk_K_r_365

   PIN u2_uk_K_r_380
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 202.65 191.49 202.75 192 ;
      END
   END u2_uk_K_r_380

   PIN u2_uk_K_r_420
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 237.05 191.49 237.15 192 ;
      END
   END u2_uk_K_r_420

   PIN FE_OFN1065_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 164.8 191.745 165 192 ;
      END
   END FE_OFN1065_n_116

   PIN FE_OFN1078_n_80338
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 432.05 191.49 432.15 192 ;
      END
   END FE_OFN1078_n_80338

   PIN FE_OFN1107_n_20850
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.45 191.49 211.55 192 ;
      END
   END FE_OFN1107_n_20850

   PIN FE_OFN1113_n_21429
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 161.45 191.49 161.55 192 ;
      END
   END FE_OFN1113_n_21429

   PIN FE_OFN1151_n_14527
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.25 191.49 188.35 192 ;
      END
   END FE_OFN1151_n_14527

   PIN FE_OFN1237_n_19800
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 332.65 0 332.75 0.51 ;
      END
   END FE_OFN1237_n_19800

   PIN FE_OFN1313_n_108168
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 447.4 191.745 447.6 192 ;
      END
   END FE_OFN1313_n_108168

   PIN FE_OFN1328_n_82601
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 110.95 0.51 111.05 ;
      END
   END FE_OFN1328_n_82601

   PIN FE_OFN15_n_106405
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.45 0 308.55 0.51 ;
      END
   END FE_OFN15_n_106405

   PIN FE_OFN1820_n_13272
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.45 191.49 79.55 192 ;
      END
   END FE_OFN1820_n_13272

   PIN FE_OFN1913_n_78988
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.25 191.49 163.35 192 ;
      END
   END FE_OFN1913_n_78988

   PIN FE_OFN217_n_15153
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 218.65 191.49 218.75 192 ;
      END
   END FE_OFN217_n_15153

   PIN FE_OFN2233_n_75724
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.25 191.49 57.35 192 ;
      END
   END FE_OFN2233_n_75724

   PIN FE_OFN2249_n_82961
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 241.25 191.49 241.35 192 ;
      END
   END FE_OFN2249_n_82961

   PIN FE_OFN2252_n_80982
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.45 191.49 188.55 192 ;
      END
   END FE_OFN2252_n_80982

   PIN FE_OFN244_n_79557
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.05 191.49 188.15 192 ;
      END
   END FE_OFN244_n_79557

   PIN FE_OFN249_n_79888
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.45 191.49 103.55 192 ;
      END
   END FE_OFN249_n_79888

   PIN FE_OFN2516_n_15149
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 308.65 191.49 308.75 192 ;
      END
   END FE_OFN2516_n_15149

   PIN FE_OFN255_n_80260
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.65 191.49 284.75 192 ;
      END
   END FE_OFN255_n_80260

   PIN FE_OFN257_n_79862
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.65 191.49 271.75 192 ;
      END
   END FE_OFN257_n_79862

   PIN FE_OFN273_n_75824
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.85 191.49 56.95 192 ;
      END
   END FE_OFN273_n_75824

   PIN FE_OFN2762_n_107068
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 452.25 191.49 452.35 192 ;
      END
   END FE_OFN2762_n_107068

   PIN FE_OFN2801_n_104989
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.55 0.51 96.65 ;
      END
   END FE_OFN2801_n_104989

   PIN FE_OFN2803_n_118632
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 376.8 191.745 377 192 ;
      END
   END FE_OFN2803_n_118632

   PIN FE_OFN3160_n_104975
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 27.25 191.49 27.35 192 ;
      END
   END FE_OFN3160_n_104975

   PIN FE_OFN3253_n_39
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 164.4 191.745 164.6 192 ;
      END
   END FE_OFN3253_n_39

   PIN FE_OFN3491_n_83012
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 213.85 191.49 213.95 192 ;
      END
   END FE_OFN3491_n_83012

   PIN FE_OFN3495_n_75992
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.85 191.49 151.95 192 ;
      END
   END FE_OFN3495_n_75992

   PIN FE_OFN3544_n_105148
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 126.85 191.49 126.95 192 ;
      END
   END FE_OFN3544_n_105148

   PIN FE_OFN3551_n_81000
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.65 191.49 185.75 192 ;
      END
   END FE_OFN3551_n_81000

   PIN FE_OFN3553_n_108480
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 490.05 191.49 490.15 192 ;
      END
   END FE_OFN3553_n_108480

   PIN FE_OFN4399_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 97.4 191.745 97.6 192 ;
      END
   END FE_OFN4399_decrypt

   PIN FE_OFN4400_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 216.8 191.745 217 192 ;
      END
   END FE_OFN4400_decrypt

   PIN FE_OFN821_n_20858
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 122.25 191.49 122.35 192 ;
      END
   END FE_OFN821_n_20858

   PIN FE_OFN865_n_15132
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 312.45 191.49 312.55 192 ;
      END
   END FE_OFN865_n_15132

   PIN g191933_p1
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 70.15 0.51 70.25 ;
      END
   END g191933_p1

   PIN g192018_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 518.05 191.49 518.15 192 ;
      END
   END g192018_da

   PIN g192018_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 518.25 191.49 518.35 192 ;
      END
   END g192018_db

   PIN g193190_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 391.65 191.49 391.75 192 ;
      END
   END g193190_p

   PIN g194055_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 452.05 191.49 452.15 192 ;
      END
   END g194055_da

   PIN g194055_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 452.05 191.49 452.15 192 ;
      END
   END g194055_db

   PIN g194626_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 249.45 191.49 249.55 192 ;
      END
   END g194626_p

   PIN g197833_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 344.45 0 344.55 0.51 ;
      END
   END g197833_da

   PIN g198664_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 227.25 191.49 227.35 192 ;
      END
   END g198664_p

   PIN g215918_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 218.05 191.49 218.15 192 ;
      END
   END g215918_p

   PIN g216302_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 215.65 191.49 215.75 192 ;
      END
   END g216302_db

   PIN g216302_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.65 191.49 198.75 192 ;
      END
   END g216302_sb

   PIN g216515_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.85 191.49 306.95 192 ;
      END
   END g216515_da

   PIN g216515_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 307.05 191.49 307.15 192 ;
      END
   END g216515_db

   PIN g216746_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 247.85 191.49 247.95 192 ;
      END
   END g216746_sb

   PIN g217136_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 73.85 191.49 73.95 192 ;
      END
   END g217136_p

   PIN g217299_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 260.45 191.49 260.55 192 ;
      END
   END g217299_p

   PIN g218012_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.45 0 44.55 0.51 ;
      END
   END g218012_p

   PIN g219309_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.25 191.49 127.35 192 ;
      END
   END g219309_p

   PIN g219396_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 295.85 191.49 295.95 192 ;
      END
   END g219396_p

   PIN g219482_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.25 191.49 104.35 192 ;
      END
   END g219482_p

   PIN g219847_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 128.05 191.49 128.15 192 ;
      END
   END g219847_p

   PIN g220720_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 357.25 191.49 357.35 192 ;
      END
   END g220720_da

   PIN g220720_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.65 191.49 79.75 192 ;
      END
   END g220720_db

   PIN g220874_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 71.05 191.49 71.15 192 ;
      END
   END g220874_db

   PIN g220874_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 63.25 191.49 63.35 192 ;
      END
   END g220874_sb

   PIN g222231_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.85 191.49 56.95 192 ;
      END
   END g222231_p

   PIN g222770_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.65 191.49 67.75 192 ;
      END
   END g222770_db

   PIN g222770_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 51.85 191.49 51.95 192 ;
      END
   END g222770_sb

   PIN g223067_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.25 191.49 81.35 192 ;
      END
   END g223067_da

   PIN g223067_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.45 191.49 81.55 192 ;
      END
   END g223067_db

   PIN g223067_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.25 191.49 80.35 192 ;
      END
   END g223067_sb

   PIN g223077_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 110.05 191.49 110.15 192 ;
      END
   END g223077_db

   PIN g223077_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.05 191.49 116.15 192 ;
      END
   END g223077_sb

   PIN g224248_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 50.65 191.49 50.75 192 ;
      END
   END g224248_db

   PIN g288145_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.85 191.49 175.95 192 ;
      END
   END g288145_p

   PIN g288651_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 85.45 191.49 85.55 192 ;
      END
   END g288651_p

   PIN g322456_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.65 191.49 140.75 192 ;
      END
   END g322456_sb

   PIN g322683_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 452.85 191.49 452.95 192 ;
      END
   END g322683_da

   PIN g322683_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 452.65 191.49 452.75 192 ;
      END
   END g322683_db

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.85 191.49 128.95 192 ;
      END
   END ispd_clk

   PIN key_c_r_30__2103
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.05 191.49 221.15 192 ;
      END
   END key_c_r_30__2103

   PIN key_c_r_32__2208
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.05 0 282.15 0.51 ;
      END
   END key_c_r_32__2208

   PIN key_c_r_32__2214
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 236.25 191.49 236.35 192 ;
      END
   END key_c_r_32__2214

   PIN key_c_r_32__2243
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 248.05 191.49 248.15 192 ;
      END
   END key_c_r_32__2243

   PIN key_c_r_33__30_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 139.15 0.51 139.25 ;
      END
   END key_c_r_33__30_

   PIN n_100299
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.65 191.49 233.75 192 ;
      END
   END n_100299

   PIN n_100477
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 283.05 191.49 283.15 192 ;
      END
   END n_100477

   PIN n_100495
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 259.45 191.49 259.55 192 ;
      END
   END n_100495

   PIN n_100662
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 241.25 191.49 241.35 192 ;
      END
   END n_100662

   PIN n_100714
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.45 191.49 260.55 192 ;
      END
   END n_100714

   PIN n_100761
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.45 191.49 282.55 192 ;
      END
   END n_100761

   PIN n_100762
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 281.85 191.49 281.95 192 ;
      END
   END n_100762

   PIN n_101445
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 390.85 191.49 390.95 192 ;
      END
   END n_101445

   PIN n_101500
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 428.05 191.49 428.15 192 ;
      END
   END n_101500

   PIN n_101504
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 402.85 191.49 402.95 192 ;
      END
   END n_101504

   PIN n_101636
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 391.05 191.49 391.15 192 ;
      END
   END n_101636

   PIN n_101645
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 410.65 191.49 410.75 192 ;
      END
   END n_101645

   PIN n_101699
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 440.05 191.49 440.15 192 ;
      END
   END n_101699

   PIN n_101768
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 400.65 191.49 400.75 192 ;
      END
   END n_101768

   PIN n_101913
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 383.05 191.49 383.15 192 ;
      END
   END n_101913

   PIN n_102201
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 440.45 191.49 440.55 192 ;
      END
   END n_102201

   PIN n_102880
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 488.65 191.49 488.75 192 ;
      END
   END n_102880

   PIN n_102908
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 199.85 191.49 199.95 192 ;
      END
   END n_102908

   PIN n_102997
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.85 191.49 248.95 192 ;
      END
   END n_102997

   PIN n_103008
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.25 0 140.35 0.51 ;
      END
   END n_103008

   PIN n_103115
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.45 191.49 152.55 192 ;
      END
   END n_103115

   PIN n_103266
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.45 191.49 284.55 192 ;
      END
   END n_103266

   PIN n_103664
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.85 191.49 282.95 192 ;
      END
   END n_103664

   PIN n_103670
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.25 191.49 260.35 192 ;
      END
   END n_103670

   PIN n_103671
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.45 191.49 271.55 192 ;
      END
   END n_103671

   PIN n_103694
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 275.05 191.49 275.15 192 ;
      END
   END n_103694

   PIN n_103802
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.65 191.49 255.75 192 ;
      END
   END n_103802

   PIN n_103837
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.25 191.49 271.35 192 ;
      END
   END n_103837

   PIN n_103855
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.85 191.49 281.95 192 ;
      END
   END n_103855

   PIN n_103882
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 253.85 191.49 253.95 192 ;
      END
   END n_103882

   PIN n_103972
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 259.45 191.49 259.55 192 ;
      END
   END n_103972

   PIN n_103998
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.05 191.49 271.15 192 ;
      END
   END n_103998

   PIN n_104090
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.05 191.49 266.15 192 ;
      END
   END n_104090

   PIN n_104111
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.85 191.49 266.95 192 ;
      END
   END n_104111

   PIN n_104147
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 282.85 191.49 282.95 192 ;
      END
   END n_104147

   PIN n_104148
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.25 191.49 245.35 192 ;
      END
   END n_104148

   PIN n_104284
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.85 191.49 270.95 192 ;
      END
   END n_104284

   PIN n_104373
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.05 191.49 260.15 192 ;
      END
   END n_104373

   PIN n_104411
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.65 191.49 270.75 192 ;
      END
   END n_104411

   PIN n_104493
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.65 191.49 267.75 192 ;
      END
   END n_104493

   PIN n_104505
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.25 191.49 255.35 192 ;
      END
   END n_104505

   PIN n_104520
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 259.85 191.49 259.95 192 ;
      END
   END n_104520

   PIN n_104588
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.25 191.49 266.35 192 ;
      END
   END n_104588

   PIN n_104625
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.05 191.49 245.15 192 ;
      END
   END n_104625

   PIN n_104873
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 463.85 191.49 463.95 192 ;
      END
   END n_104873

   PIN n_105003
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 228.45 191.49 228.55 192 ;
      END
   END n_105003

   PIN n_105099
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 259.25 191.49 259.35 192 ;
      END
   END n_105099

   PIN n_105150
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 356.85 191.49 356.95 192 ;
      END
   END n_105150

   PIN n_105176
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.95 0.51 60.05 ;
      END
   END n_105176

   PIN n_105284
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.75 0.51 59.85 ;
      END
   END n_105284

   PIN n_105286
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.75 0.51 83.85 ;
      END
   END n_105286

   PIN n_105287
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 96.1 0.255 96.3 ;
      END
   END n_105287

   PIN n_105353
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 60.95 0.51 61.05 ;
      END
   END n_105353

   PIN n_105423
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.45 0 224.55 0.51 ;
      END
   END n_105423

   PIN n_105424
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 216.25 191.49 216.35 192 ;
      END
   END n_105424

   PIN n_105451
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.15 0.51 68.25 ;
      END
   END n_105451

   PIN n_105486
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 363.65 191.49 363.75 192 ;
      END
   END n_105486

   PIN n_105503
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.85 0 212.95 0.51 ;
      END
   END n_105503

   PIN n_105531
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 68.75 0.51 68.85 ;
      END
   END n_105531

   PIN n_105540
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.05 0 212.15 0.51 ;
      END
   END n_105540

   PIN n_105541
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.45 0 221.55 0.51 ;
      END
   END n_105541

   PIN n_105547
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.55 0.51 83.65 ;
      END
   END n_105547

   PIN n_105552
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 505.65 191.49 505.75 192 ;
      END
   END n_105552

   PIN n_105593
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 192.45 0 192.55 0.51 ;
      END
   END n_105593

   PIN n_105596
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.45 0 284.55 0.51 ;
      END
   END n_105596

   PIN n_105632
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.85 0 211.95 0.51 ;
      END
   END n_105632

   PIN n_105634
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 60.35 0.51 60.45 ;
      END
   END n_105634

   PIN n_105645
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 198.05 0 198.15 0.51 ;
      END
   END n_105645

   PIN n_105648
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 367.05 191.49 367.15 192 ;
      END
   END n_105648

   PIN n_105678
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 505.45 191.49 505.55 192 ;
      END
   END n_105678

   PIN n_105694
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 81.15 0.51 81.25 ;
      END
   END n_105694

   PIN n_105696
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 228.45 0 228.55 0.51 ;
      END
   END n_105696

   PIN n_105707
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 364.05 191.49 364.15 192 ;
      END
   END n_105707

   PIN n_105715
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 250.05 0 250.15 0.51 ;
      END
   END n_105715

   PIN n_105739
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 200.85 0 200.95 0.51 ;
      END
   END n_105739

   PIN n_105749
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.45 0 248.55 0.51 ;
      END
   END n_105749

   PIN n_105788
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 94.95 0.51 95.05 ;
      END
   END n_105788

   PIN n_105875
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 67.95 0.51 68.05 ;
      END
   END n_105875

   PIN n_105910
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.35 0.51 70.45 ;
      END
   END n_105910

   PIN n_105912
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 215.25 0 215.35 0.51 ;
      END
   END n_105912

   PIN n_105916
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.25 0 224.35 0.51 ;
      END
   END n_105916

   PIN n_105937
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 67.75 0.51 67.85 ;
      END
   END n_105937

   PIN n_105995
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 236.65 0 236.75 0.51 ;
      END
   END n_105995

   PIN n_106012
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 392.65 191.49 392.75 192 ;
      END
   END n_106012

   PIN n_106014
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 376.05 191.49 376.15 192 ;
      END
   END n_106014

   PIN n_106037
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 81.75 0.51 81.85 ;
      END
   END n_106037

   PIN n_106057
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 392.05 191.49 392.15 192 ;
      END
   END n_106057

   PIN n_106089
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 67.55 0.51 67.65 ;
      END
   END n_106089

   PIN n_106090
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.55 0.51 59.65 ;
      END
   END n_106090

   PIN n_106099
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.35 0.51 83.45 ;
      END
   END n_106099

   PIN n_106148
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 365.65 191.49 365.75 192 ;
      END
   END n_106148

   PIN n_106153
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.35 0.51 59.45 ;
      END
   END n_106153

   PIN n_106158
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.45 0 176.55 0.51 ;
      END
   END n_106158

   PIN n_106159
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.45 0 164.55 0.51 ;
      END
   END n_106159

   PIN n_106162
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.95 0.51 71.05 ;
      END
   END n_106162

   PIN n_106163
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 67.35 0.51 67.45 ;
      END
   END n_106163

   PIN n_106166
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.75 0.51 70.85 ;
      END
   END n_106166

   PIN n_106171
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.05 0 185.15 0.51 ;
      END
   END n_106171

   PIN n_106182
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 384.65 191.49 384.75 192 ;
      END
   END n_106182

   PIN n_106184
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 502.65 191.49 502.75 192 ;
      END
   END n_106184

   PIN n_106194
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 187.85 0 187.95 0.51 ;
      END
   END n_106194

   PIN n_106196
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.75 0.51 51.85 ;
      END
   END n_106196

   PIN n_106200
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.45 0 212.55 0.51 ;
      END
   END n_106200

   PIN n_106207
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 398.65 191.49 398.75 192 ;
      END
   END n_106207

   PIN n_106208
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 379.85 191.49 379.95 192 ;
      END
   END n_106208

   PIN n_106220
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 59.15 0.51 59.25 ;
      END
   END n_106220

   PIN n_106224
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.25 0 152.35 0.51 ;
      END
   END n_106224

   PIN n_106247
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 384.25 191.49 384.35 192 ;
      END
   END n_106247

   PIN n_106253
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 60.75 0.51 60.85 ;
      END
   END n_106253

   PIN n_106258
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.55 0.51 70.65 ;
      END
   END n_106258

   PIN n_106273
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 60.55 0.51 60.65 ;
      END
   END n_106273

   PIN n_106306
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 391.45 191.49 391.55 192 ;
      END
   END n_106306

   PIN n_106327
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.55 0.51 71.65 ;
      END
   END n_106327

   PIN n_106329
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.95 0.51 84.05 ;
      END
   END n_106329

   PIN n_106337
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 60.15 0.51 60.25 ;
      END
   END n_106337

   PIN n_106361
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 201.45 0 201.55 0.51 ;
      END
   END n_106361

   PIN n_106445
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 206.45 0 206.55 0.51 ;
      END
   END n_106445

   PIN n_106450
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.85 0 199.95 0.51 ;
      END
   END n_106450

   PIN n_106452
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.95 0.51 59.05 ;
      END
   END n_106452

   PIN n_106488
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 384.05 191.49 384.15 192 ;
      END
   END n_106488

   PIN n_106510
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 373.45 191.49 373.55 192 ;
      END
   END n_106510

   PIN n_106526
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 67.15 0.51 67.25 ;
      END
   END n_106526

   PIN n_106531
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 143.65 0 143.75 0.51 ;
      END
   END n_106531

   PIN n_106533
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 392.45 191.49 392.55 192 ;
      END
   END n_106533

   PIN n_106568
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.25 0 176.35 0.51 ;
      END
   END n_106568

   PIN n_106586
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 183.65 0 183.75 0.51 ;
      END
   END n_106586

   PIN n_106596
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.65 0 272.75 0.51 ;
      END
   END n_106596

   PIN n_106597
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.25 0 164.35 0.51 ;
      END
   END n_106597

   PIN n_106601
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 160.65 0 160.75 0.51 ;
      END
   END n_106601

   PIN n_106603
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 7.15 0.51 7.25 ;
      END
   END n_106603

   PIN n_106608
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.65 0 199.75 0.51 ;
      END
   END n_106608

   PIN n_106629
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 379.65 191.49 379.75 192 ;
      END
   END n_106629

   PIN n_106649
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.75 0.51 58.85 ;
      END
   END n_106649

   PIN n_106661
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 373.65 191.49 373.75 192 ;
      END
   END n_106661

   PIN n_106663
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 236.45 0 236.55 0.51 ;
      END
   END n_106663

   PIN n_106710
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 392.25 191.49 392.35 192 ;
      END
   END n_106710

   PIN n_106714
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.95 0.51 39.05 ;
      END
   END n_106714

   PIN n_106751
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 379.45 191.49 379.55 192 ;
      END
   END n_106751

   PIN n_106817
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.65 0 140.75 0.51 ;
      END
   END n_106817

   PIN n_106818
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 488.85 191.49 488.95 192 ;
      END
   END n_106818

   PIN n_106840
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.45 0 140.55 0.51 ;
      END
   END n_106840

   PIN n_106900
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 501.05 191.49 501.15 192 ;
      END
   END n_106900

   PIN n_107024
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 517.05 191.49 517.15 192 ;
      END
   END n_107024

   PIN n_107054
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 51.15 523 51.25 ;
      END
   END n_107054

   PIN n_107067
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 486.65 191.49 486.75 192 ;
      END
   END n_107067

   PIN n_107081
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 501.65 191.49 501.75 192 ;
      END
   END n_107081

   PIN n_107097
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 502.85 191.49 502.95 192 ;
      END
   END n_107097

   PIN n_107129
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 472.25 191.49 472.35 192 ;
      END
   END n_107129

   PIN n_107136
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 475.25 191.49 475.35 192 ;
      END
   END n_107136

   PIN n_107146
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 487.45 191.49 487.55 192 ;
      END
   END n_107146

   PIN n_107190
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 467.8 191.745 468 192 ;
      END
   END n_107190

   PIN n_107250
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 501.25 191.49 501.35 192 ;
      END
   END n_107250

   PIN n_107253
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 502.05 191.49 502.15 192 ;
      END
   END n_107253

   PIN n_107341
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 502.25 191.49 502.35 192 ;
      END
   END n_107341

   PIN n_107345
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 509.85 0 509.95 0.51 ;
      END
   END n_107345

   PIN n_107369
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 140.95 523 141.05 ;
      END
   END n_107369

   PIN n_107412
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 502.45 191.49 502.55 192 ;
      END
   END n_107412

   PIN n_107462
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 124.95 523 125.05 ;
      END
   END n_107462

   PIN n_107486
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 139.15 523 139.25 ;
      END
   END n_107486

   PIN n_107495
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 514.05 191.49 514.15 192 ;
      END
   END n_107495

   PIN n_107519
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 95.15 523 95.25 ;
      END
   END n_107519

   PIN n_107577
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 440.65 0 440.75 0.51 ;
      END
   END n_107577

   PIN n_107602
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 501.45 191.49 501.55 192 ;
      END
   END n_107602

   PIN n_107611
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 487.45 191.49 487.55 192 ;
      END
   END n_107611

   PIN n_107634
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 465.85 0 465.95 0.51 ;
      END
   END n_107634

   PIN n_107640
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 502.65 191.49 502.75 192 ;
      END
   END n_107640

   PIN n_107641
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 138.95 523 139.05 ;
      END
   END n_107641

   PIN n_107652
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 500.85 191.49 500.95 192 ;
      END
   END n_107652

   PIN n_107656
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 71.95 523 72.05 ;
      END
   END n_107656

   PIN n_107660
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 497.25 191.49 497.35 192 ;
      END
   END n_107660

   PIN n_107674
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 168.95 523 169.05 ;
      END
   END n_107674

   PIN n_107677
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.745 110.9 523 111.1 ;
      END
   END n_107677

   PIN n_107723
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 463.65 191.49 463.75 192 ;
      END
   END n_107723

   PIN n_107738
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 512.25 0 512.35 0.51 ;
      END
   END n_107738

   PIN n_107746
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 464.65 191.49 464.75 192 ;
      END
   END n_107746

   PIN n_107782
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 487.65 191.49 487.75 192 ;
      END
   END n_107782

   PIN n_107829
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 356.45 0 356.55 0.51 ;
      END
   END n_107829

   PIN n_107928
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 487.85 191.49 487.95 192 ;
      END
   END n_107928

   PIN n_107943
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 22.95 523 23.05 ;
      END
   END n_107943

   PIN n_107996
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 83.75 523 83.85 ;
      END
   END n_107996

   PIN n_108012
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 501.25 191.49 501.35 192 ;
      END
   END n_108012

   PIN n_108045
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 35.95 523 36.05 ;
      END
   END n_108045

   PIN n_108049
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 493.65 191.49 493.75 192 ;
      END
   END n_108049

   PIN n_108137
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 488.25 191.49 488.35 192 ;
      END
   END n_108137

   PIN n_108148
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 479.45 191.49 479.55 192 ;
      END
   END n_108148

   PIN n_108191
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 464.05 191.49 464.15 192 ;
      END
   END n_108191

   PIN n_108245
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 488.45 0 488.55 0.51 ;
      END
   END n_108245

   PIN n_108254
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 451.85 191.49 451.95 192 ;
      END
   END n_108254

   PIN n_108278
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 483.05 191.49 483.15 192 ;
      END
   END n_108278

   PIN n_108295
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 71.75 523 71.85 ;
      END
   END n_108295

   PIN n_108407
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 81.15 523 81.25 ;
      END
   END n_108407

   PIN n_108410
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 522.49 94.95 523 95.05 ;
      END
   END n_108410

   PIN n_108418
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 464.25 191.49 464.35 192 ;
      END
   END n_108418

   PIN n_108449
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 464.85 191.49 464.95 192 ;
      END
   END n_108449

   PIN n_108499
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 493.05 191.49 493.15 192 ;
      END
   END n_108499

   PIN n_109142
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.45 191.49 116.55 192 ;
      END
   END n_109142

   PIN n_109209
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 111.85 191.49 111.95 192 ;
      END
   END n_109209

   PIN n_116820
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 400.85 191.49 400.95 192 ;
      END
   END n_116820

   PIN n_117788
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 189.25 191.49 189.35 192 ;
      END
   END n_117788

   PIN n_118032
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 513.85 191.49 513.95 192 ;
      END
   END n_118032

   PIN n_118355
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.85 191.49 292.95 192 ;
      END
   END n_118355

   PIN n_118357
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 275.25 191.49 275.35 192 ;
      END
   END n_118357

   PIN n_118359
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.45 191.49 272.55 192 ;
      END
   END n_118359

   PIN n_118364
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 296.65 191.49 296.75 192 ;
      END
   END n_118364

   PIN n_118371
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.65 191.49 285.75 192 ;
      END
   END n_118371

   PIN n_118636
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 391.85 191.49 391.95 192 ;
      END
   END n_118636

   PIN n_118642
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 367.85 191.49 367.95 192 ;
      END
   END n_118642

   PIN n_118707
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 308.45 191.49 308.55 192 ;
      END
   END n_118707

   PIN n_126097
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 412.85 191.49 412.95 192 ;
      END
   END n_126097

   PIN n_13376
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 96.05 191.49 96.15 192 ;
      END
   END n_13376

   PIN n_13380
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.25 191.49 124.35 192 ;
      END
   END n_13380

   PIN n_13382
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 145.45 191.49 145.55 192 ;
      END
   END n_13382

   PIN n_13477
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.65 191.49 139.75 192 ;
      END
   END n_13477

   PIN n_13479
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 139.65 191.49 139.75 192 ;
      END
   END n_13479

   PIN n_13482
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.45 191.49 139.55 192 ;
      END
   END n_13482

   PIN n_13488
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 109.45 191.49 109.55 192 ;
      END
   END n_13488

   PIN n_13521
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 3.05 191.49 3.15 192 ;
      END
   END n_13521

   PIN n_13606
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 127.25 191.49 127.35 192 ;
      END
   END n_13606

   PIN n_13710
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 217.85 191.49 217.95 192 ;
      END
   END n_13710

   PIN n_137147
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.55 0.51 38.65 ;
      END
   END n_137147

   PIN n_137154
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.65 191.49 20.75 192 ;
      END
   END n_137154

   PIN n_13741
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.85 191.49 115.95 192 ;
      END
   END n_13741

   PIN n_13754
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 110.25 191.49 110.35 192 ;
      END
   END n_13754

   PIN n_13841
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 204.25 191.49 204.35 192 ;
      END
   END n_13841

   PIN n_13861
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 128.25 191.49 128.35 192 ;
      END
   END n_13861

   PIN n_13872
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 222.05 191.49 222.15 192 ;
      END
   END n_13872

   PIN n_13981
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.65 191.49 177.75 192 ;
      END
   END n_13981

   PIN n_14011
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 185.85 191.49 185.95 192 ;
      END
   END n_14011

   PIN n_14014
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.05 191.49 177.15 192 ;
      END
   END n_14014

   PIN n_14026
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 151.65 191.49 151.75 192 ;
      END
   END n_14026

   PIN n_14129
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 132.25 191.49 132.35 192 ;
      END
   END n_14129

   PIN n_14373
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 127.45 191.49 127.55 192 ;
      END
   END n_14373

   PIN n_14379
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 150.85 191.49 150.95 192 ;
      END
   END n_14379

   PIN n_14517
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 179.65 191.49 179.75 192 ;
      END
   END n_14517

   PIN n_14520
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 162.25 191.49 162.35 192 ;
      END
   END n_14520

   PIN n_14525
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 166.65 191.49 166.75 192 ;
      END
   END n_14525

   PIN n_15151
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.45 191.49 164.55 192 ;
      END
   END n_15151

   PIN n_15369
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.05 191.49 212.15 192 ;
      END
   END n_15369

   PIN n_212521
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 160.25 191.49 160.35 192 ;
      END
   END n_212521

   PIN n_21351
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.45 191.49 57.55 192 ;
      END
   END n_21351

   PIN n_21398
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.65 191.49 188.75 192 ;
      END
   END n_21398

   PIN n_21430
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.85 191.49 164.95 192 ;
      END
   END n_21430

   PIN n_75475
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 85.05 191.49 85.15 192 ;
      END
   END n_75475

   PIN n_75713
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 96.85 191.49 96.95 192 ;
      END
   END n_75713

   PIN n_75715
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 85.25 191.49 85.35 192 ;
      END
   END n_75715

   PIN n_75770
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 192.25 191.49 192.35 192 ;
      END
   END n_75770

   PIN n_75788
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 153.45 191.49 153.55 192 ;
      END
   END n_75788

   PIN n_76012
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 15.85 191.49 15.95 192 ;
      END
   END n_76012

   PIN n_76214
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 29.2 191.745 29.4 192 ;
      END
   END n_76214

   PIN n_76298
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.45 191.49 44.55 192 ;
      END
   END n_76298

   PIN n_76529
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 67.25 191.49 67.35 192 ;
      END
   END n_76529

   PIN n_76816
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 45.05 191.49 45.15 192 ;
      END
   END n_76816

   PIN n_76865
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.05 191.49 10.15 192 ;
      END
   END n_76865

   PIN n_76896
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 58.05 191.49 58.15 192 ;
      END
   END n_76896

   PIN n_76931
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 57.05 191.49 57.15 192 ;
      END
   END n_76931

   PIN n_76932
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 53.25 191.49 53.35 192 ;
      END
   END n_76932

   PIN n_76935
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 67.45 191.49 67.55 192 ;
      END
   END n_76935

   PIN n_77062
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 53.45 191.49 53.55 192 ;
      END
   END n_77062

   PIN n_77148
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 43.85 191.49 43.95 192 ;
      END
   END n_77148

   PIN n_77280
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 23.25 191.49 23.35 192 ;
      END
   END n_77280

   PIN n_77331
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 57.85 191.49 57.95 192 ;
      END
   END n_77331

   PIN n_77392
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44 191.745 44.2 192 ;
      END
   END n_77392

   PIN n_77415
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 3.25 191.49 3.35 192 ;
      END
   END n_77415

   PIN n_77416
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44.45 191.49 44.55 192 ;
      END
   END n_77416

   PIN n_77722
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.85 191.49 31.95 192 ;
      END
   END n_77722

   PIN n_77723
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.45 191.49 40.55 192 ;
      END
   END n_77723

   PIN n_77759
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 44.65 191.49 44.75 192 ;
      END
   END n_77759

   PIN n_77771
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.05 191.49 44.15 192 ;
      END
   END n_77771

   PIN n_77821
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 32.25 191.49 32.35 192 ;
      END
   END n_77821

   PIN n_77947
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 16.05 191.49 16.15 192 ;
      END
   END n_77947

   PIN n_78815
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.85 191.49 20.95 192 ;
      END
   END n_78815

   PIN n_78831
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 164.05 191.49 164.15 192 ;
      END
   END n_78831

   PIN n_78876
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 297.05 191.49 297.15 192 ;
      END
   END n_78876

   PIN n_78916
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 223.85 191.49 223.95 192 ;
      END
   END n_78916

   PIN n_78927
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.65 191.49 115.75 192 ;
      END
   END n_78927

   PIN n_78965
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 169.65 191.49 169.75 192 ;
      END
   END n_78965

   PIN n_78977
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.25 191.49 285.35 192 ;
      END
   END n_78977

   PIN n_78990
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 177.45 191.49 177.55 192 ;
      END
   END n_78990

   PIN n_78998
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.85 191.49 163.95 192 ;
      END
   END n_78998

   PIN n_79103
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 160.45 191.49 160.55 192 ;
      END
   END n_79103

   PIN n_79120
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.45 191.49 128.55 192 ;
      END
   END n_79120

   PIN n_79137
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.05 191.49 285.15 192 ;
      END
   END n_79137

   PIN n_79146
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.85 191.49 188.95 192 ;
      END
   END n_79146

   PIN n_79180
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 344.65 191.49 344.75 192 ;
      END
   END n_79180

   PIN n_79289
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 425.25 191.49 425.35 192 ;
      END
   END n_79289

   PIN n_79305
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.85 191.49 127.95 192 ;
      END
   END n_79305

   PIN n_79354
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 224.25 191.49 224.35 192 ;
      END
   END n_79354

   PIN n_79364
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.05 191.49 272.15 192 ;
      END
   END n_79364

   PIN n_79384
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 324.05 191.49 324.15 192 ;
      END
   END n_79384

   PIN n_79386
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 144.05 191.49 144.15 192 ;
      END
   END n_79386

   PIN n_79389
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 184.05 191.49 184.15 192 ;
      END
   END n_79389

   PIN n_79393
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 89.25 191.49 89.35 192 ;
      END
   END n_79393

   PIN n_79422
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 290.65 191.49 290.75 192 ;
      END
   END n_79422

   PIN n_79423
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 238.05 191.49 238.15 192 ;
      END
   END n_79423

   PIN n_79461
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 432.25 191.49 432.35 192 ;
      END
   END n_79461

   PIN n_79469
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 156.85 191.49 156.95 192 ;
      END
   END n_79469

   PIN n_79525
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.45 191.49 285.55 192 ;
      END
   END n_79525

   PIN n_79565
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 349.45 0 349.55 0.51 ;
      END
   END n_79565

   PIN n_79566
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 271.85 191.49 271.95 192 ;
      END
   END n_79566

   PIN n_79570
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 89.65 191.49 89.75 192 ;
      END
   END n_79570

   PIN n_79571
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 126.65 191.49 126.75 192 ;
      END
   END n_79571

   PIN n_79575
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 404.25 191.49 404.35 192 ;
      END
   END n_79575

   PIN n_79576
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 128.45 191.49 128.55 192 ;
      END
   END n_79576

   PIN n_79622
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.25 191.49 272.35 192 ;
      END
   END n_79622

   PIN n_79636
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.45 191.49 248.55 192 ;
      END
   END n_79636

   PIN n_79679
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 248.25 191.49 248.35 192 ;
      END
   END n_79679

   PIN n_79720
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 324.45 191.49 324.55 192 ;
      END
   END n_79720

   PIN n_79734
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.85 191.49 283.95 192 ;
      END
   END n_79734

   PIN n_79739
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 284.25 191.49 284.35 192 ;
      END
   END n_79739

   PIN n_79776
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 436.65 191.49 436.75 192 ;
      END
   END n_79776

   PIN n_79781
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 401.65 191.49 401.75 192 ;
      END
   END n_79781

   PIN n_79802
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 237.25 191.49 237.35 192 ;
      END
   END n_79802

   PIN n_79857
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.25 191.49 105.35 192 ;
      END
   END n_79857

   PIN n_79870
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.45 191.49 104.55 192 ;
      END
   END n_79870

   PIN n_79886
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 117.85 191.49 117.95 192 ;
      END
   END n_79886

   PIN n_79924
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 415.45 191.49 415.55 192 ;
      END
   END n_79924

   PIN n_79933
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 429.25 191.49 429.35 192 ;
      END
   END n_79933

   PIN n_79945
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 302.05 191.49 302.15 192 ;
      END
   END n_79945

   PIN n_79963
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 247.25 191.49 247.35 192 ;
      END
   END n_79963

   PIN n_79967
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.65 191.49 116.75 192 ;
      END
   END n_79967

   PIN n_80003
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 344.85 191.49 344.95 192 ;
      END
   END n_80003

   PIN n_80022
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 136.65 191.49 136.75 192 ;
      END
   END n_80022

   PIN n_80032
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 211.85 191.49 211.95 192 ;
      END
   END n_80032

   PIN n_80060
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 445.85 191.49 445.95 192 ;
      END
   END n_80060

   PIN n_80067
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 416.85 191.49 416.95 192 ;
      END
   END n_80067

   PIN n_80068
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 417.85 191.49 417.95 192 ;
      END
   END n_80068

   PIN n_80096
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 424.45 191.49 424.55 192 ;
      END
   END n_80096

   PIN n_80115
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.05 191.49 284.15 192 ;
      END
   END n_80115

   PIN n_80137
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 337.65 191.49 337.75 192 ;
      END
   END n_80137

   PIN n_80149
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.45 191.49 212.55 192 ;
      END
   END n_80149

   PIN n_80206
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 408 191.745 408.2 192 ;
      END
   END n_80206

   PIN n_80245
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 415.25 191.49 415.35 192 ;
      END
   END n_80245

   PIN n_80249
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.05 191.49 128.15 192 ;
      END
   END n_80249

   PIN n_80253
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.85 191.49 140.95 192 ;
      END
   END n_80253

   PIN n_80274
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 440.25 191.49 440.35 192 ;
      END
   END n_80274

   PIN n_80282
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 212.05 191.49 212.15 192 ;
      END
   END n_80282

   PIN n_80325
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 427.25 191.49 427.35 192 ;
      END
   END n_80325

   PIN n_80329
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 416.65 191.49 416.75 192 ;
      END
   END n_80329

   PIN n_80387
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 284.05 191.49 284.15 192 ;
      END
   END n_80387

   PIN n_80393
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 265.45 191.49 265.55 192 ;
      END
   END n_80393

   PIN n_80399
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 314.05 191.49 314.15 192 ;
      END
   END n_80399

   PIN n_80401
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 142.65 191.49 142.75 192 ;
      END
   END n_80401

   PIN n_80404
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 104.65 191.49 104.75 192 ;
      END
   END n_80404

   PIN n_80408
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 403.65 191.49 403.75 192 ;
      END
   END n_80408

   PIN n_80412
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 416.45 191.49 416.55 192 ;
      END
   END n_80412

   PIN n_80425
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 263.65 191.49 263.75 192 ;
      END
   END n_80425

   PIN n_80429
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 427.65 191.49 427.75 192 ;
      END
   END n_80429

   PIN n_80504
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 222.65 191.49 222.75 192 ;
      END
   END n_80504

   PIN n_80520
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 116.85 191.49 116.95 192 ;
      END
   END n_80520

   PIN n_80538
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 424.25 191.49 424.35 192 ;
      END
   END n_80538

   PIN n_80551
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 200.85 191.49 200.95 192 ;
      END
   END n_80551

   PIN n_80557
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 186.45 191.49 186.55 192 ;
      END
   END n_80557

   PIN n_80619
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 79.45 191.49 79.55 192 ;
      END
   END n_80619

   PIN n_80631
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 280.45 191.49 280.55 192 ;
      END
   END n_80631

   PIN n_80640
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 408.25 191.49 408.35 192 ;
      END
   END n_80640

   PIN n_80682
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 309.85 191.49 309.95 192 ;
      END
   END n_80682

   PIN n_80694
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.05 191.49 176.15 192 ;
      END
   END n_80694

   PIN n_80734
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 141.05 191.49 141.15 192 ;
      END
   END n_80734

   PIN n_80743
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.25 191.49 282.35 192 ;
      END
   END n_80743

   PIN n_80759
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 156.05 191.49 156.15 192 ;
      END
   END n_80759

   PIN n_80763
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 229.25 191.49 229.35 192 ;
      END
   END n_80763

   PIN n_80777
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 419.85 191.49 419.95 192 ;
      END
   END n_80777

   PIN n_80788
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.25 0 260.35 0.51 ;
      END
   END n_80788

   PIN n_80817
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 357.05 191.49 357.15 192 ;
      END
   END n_80817

   PIN n_80905
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.25 191.49 176.35 192 ;
      END
   END n_80905

   PIN n_80956
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 152.25 191.49 152.35 192 ;
      END
   END n_80956

   PIN n_81032
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 238.65 191.49 238.75 192 ;
      END
   END n_81032

   PIN n_81118
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285 191.745 285.2 192 ;
      END
   END n_81118

   PIN n_81188
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 296.85 191.49 296.95 192 ;
      END
   END n_81188

   PIN n_81261
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 296.25 191.49 296.35 192 ;
      END
   END n_81261

   PIN n_81264
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.15 0.51 38.25 ;
      END
   END n_81264

   PIN n_81273
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 44.05 0 44.15 0.51 ;
      END
   END n_81273

   PIN n_81298
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 72.25 191.49 72.35 192 ;
      END
   END n_81298

   PIN n_81301
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 310.85 191.49 310.95 192 ;
      END
   END n_81301

   PIN n_81360
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.05 191.49 55.15 192 ;
      END
   END n_81360

   PIN n_81395
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.85 191.49 284.95 192 ;
      END
   END n_81395

   PIN n_81420
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.3 0.255 23.5 ;
      END
   END n_81420

   PIN n_81431
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 22.35 0.51 22.45 ;
      END
   END n_81431

   PIN n_81462
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 58.55 0.51 58.65 ;
      END
   END n_81462

   PIN n_81477
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 284.45 191.49 284.55 192 ;
      END
   END n_81477

   PIN n_81478
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 284.25 191.49 284.35 192 ;
      END
   END n_81478

   PIN n_81503
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.95 0.51 38.05 ;
      END
   END n_81503

   PIN n_81504
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 23.75 0.51 23.85 ;
      END
   END n_81504

   PIN n_81590
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 229.05 191.49 229.15 192 ;
      END
   END n_81590

   PIN n_81626
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 38.75 0.51 38.85 ;
      END
   END n_81626

   PIN n_81646
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 342.85 191.49 342.95 192 ;
      END
   END n_81646

   PIN n_81668
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 6.95 0.51 7.05 ;
      END
   END n_81668

   PIN n_81761
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.15 0.51 25.25 ;
      END
   END n_81761

   PIN n_81776
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 237.65 191.49 237.75 192 ;
      END
   END n_81776

   PIN n_81799
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.75 0.51 37.85 ;
      END
   END n_81799

   PIN n_81886
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285.65 191.49 285.75 192 ;
      END
   END n_81886

   PIN n_81905
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 306.25 191.49 306.35 192 ;
      END
   END n_81905

   PIN n_81907
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 295.65 191.49 295.75 192 ;
      END
   END n_81907

   PIN n_81908
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 295.45 191.49 295.55 192 ;
      END
   END n_81908

   PIN n_81955
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.95 0.51 25.05 ;
      END
   END n_81955

   PIN n_82085
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 317.85 191.49 317.95 192 ;
      END
   END n_82085

   PIN n_82109
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.55 0.51 24.65 ;
      END
   END n_82109

   PIN n_82147
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.55 0.51 37.65 ;
      END
   END n_82147

   PIN n_82168
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.55 0.51 51.65 ;
      END
   END n_82168

   PIN n_82173
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 325.05 191.49 325.15 192 ;
      END
   END n_82173

   PIN n_82174
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 242.25 191.49 242.35 192 ;
      END
   END n_82174

   PIN n_82178
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.65 191.49 283.75 192 ;
      END
   END n_82178

   PIN n_82215
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.35 0.51 51.45 ;
      END
   END n_82215

   PIN n_82244
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 260.85 191.49 260.95 192 ;
      END
   END n_82244

   PIN n_82268
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 285.85 191.49 285.95 192 ;
      END
   END n_82268

   PIN n_82282
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 34.75 0.51 34.85 ;
      END
   END n_82282

   PIN n_82287
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 24.35 0.51 24.45 ;
      END
   END n_82287

   PIN n_82291
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.65 0 55.75 0.51 ;
      END
   END n_82291

   PIN n_82311
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 297.25 191.49 297.35 192 ;
      END
   END n_82311

   PIN n_82329
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 37.35 0.51 37.45 ;
      END
   END n_82329

   PIN n_82352
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 248.45 191.49 248.55 192 ;
      END
   END n_82352

   PIN n_82357
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.25 0 49.35 0.51 ;
      END
   END n_82357

   PIN n_82374
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 25.35 0.51 25.45 ;
      END
   END n_82374

   PIN n_82375
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 67.65 191.49 67.75 192 ;
      END
   END n_82375

   PIN n_82412
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 330.25 191.49 330.35 192 ;
      END
   END n_82412

   PIN n_82417
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 296.05 191.49 296.15 192 ;
      END
   END n_82417

   PIN n_82424
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 347.65 191.49 347.75 192 ;
      END
   END n_82424

   PIN n_82432
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 297.45 191.49 297.55 192 ;
      END
   END n_82432

   PIN n_82451
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 90.45 191.49 90.55 192 ;
      END
   END n_82451

   PIN n_82505
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 58.25 191.49 58.35 192 ;
      END
   END n_82505

   PIN n_82562
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 315.25 191.49 315.35 192 ;
      END
   END n_82562

   PIN n_82586
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 260.65 191.49 260.75 192 ;
      END
   END n_82586

   PIN n_82645
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 84.15 0.51 84.25 ;
      END
   END n_82645

   PIN n_82650
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 300.25 191.49 300.35 192 ;
      END
   END n_82650

   PIN n_82678
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 351.05 191.49 351.15 192 ;
      END
   END n_82678

   PIN n_82679
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 78.65 191.49 78.75 192 ;
      END
   END n_82679

   PIN n_82698
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 95.35 0.51 95.45 ;
      END
   END n_82698

   PIN n_82738
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 91.25 191.49 91.35 192 ;
      END
   END n_82738

   PIN n_82745
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.65 191.49 81.75 192 ;
      END
   END n_82745

   PIN n_82764
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 81.85 191.49 81.95 192 ;
      END
   END n_82764

   PIN n_82769
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.65 191.49 282.75 192 ;
      END
   END n_82769

   PIN n_82770
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 261.05 191.49 261.15 192 ;
      END
   END n_82770

   PIN n_83142
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 218.45 191.49 218.55 192 ;
      END
   END n_83142

   PIN n_83215
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 404.25 191.49 404.35 192 ;
      END
   END n_83215

   PIN n_84346
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 413.85 191.49 413.95 192 ;
      END
   END n_84346

   PIN n_84639
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 416.25 191.49 416.35 192 ;
      END
   END n_84639

   PIN n_84673
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 439.45 191.49 439.55 192 ;
      END
   END n_84673

   PIN n_84781
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 397.05 191.49 397.15 192 ;
      END
   END n_84781

   PIN n_84844
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 344.05 191.49 344.15 192 ;
      END
   END n_84844

   PIN n_99925
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 271.45 191.49 271.55 192 ;
      END
   END n_99925

   PIN stage2_out_3228
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 8.65 191.49 8.75 192 ;
      END
   END stage2_out_3228

   PIN stage2_out_3231
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 185.15 0.51 185.25 ;
      END
   END stage2_out_3231

   PIN stage2_out_3237
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 154.95 0.51 155.05 ;
      END
   END stage2_out_3237

   PIN stage2_out_3238
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.45 191.49 32.55 192 ;
      END
   END stage2_out_3238

   PIN stage2_out_3262
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 80.45 191.49 80.55 192 ;
      END
   END stage2_out_3262

   PIN u1_L14_20_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 138.95 0.51 139.05 ;
      END
   END u1_L14_20_

   PIN u1_R13_16_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 124.95 0.51 125.05 ;
      END
   END u1_R13_16_

   PIN u1_R13_29_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 184.95 0.51 185.05 ;
      END
   END u1_R13_29_

   PIN u1_R13_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 168.95 0.51 169.05 ;
      END
   END u1_R13_6_

   PIN u2_IP_32_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 185.35 0.51 185.45 ;
      END
   END u2_IP_32_

   PIN u2_IP_64__1271
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 100.25 191.49 100.35 192 ;
      END
   END u2_IP_64__1271

   PIN u2_IP_64__1272
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 142.85 191.49 142.95 192 ;
      END
   END u2_IP_64__1272

   PIN u2_IP_64__1273
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.85 191.49 106.95 192 ;
      END
   END u2_IP_64__1273

   PIN u2_IP_64__1278
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 56.65 191.49 56.75 192 ;
      END
   END u2_IP_64__1278

   PIN u2_IP_64__1280
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 117.25 191.49 117.35 192 ;
      END
   END u2_IP_64__1280

   PIN u2_IP_64__1282
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 10.25 191.49 10.35 192 ;
      END
   END u2_IP_64__1282

   PIN u2_IP_64__1286
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 68.25 191.49 68.35 192 ;
      END
   END u2_IP_64__1286

   PIN u2_L0_26_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.65 191.49 163.75 192 ;
      END
   END u2_L0_26_

   PIN u2_L0_31_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 188.25 191.49 188.35 192 ;
      END
   END u2_L0_31_

   PIN u2_L0_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.65 191.49 199.75 192 ;
      END
   END u2_L0_7_

   PIN u2_L0_9_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 247.05 191.49 247.15 192 ;
      END
   END u2_L0_9_

   PIN u2_L0_reg_10__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 127.65 191.49 127.75 192 ;
      END
   END u2_L0_reg_10__Q

   PIN u2_L10_27_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 224.65 191.49 224.75 192 ;
      END
   END u2_L10_27_

   PIN u2_L10_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 259.05 191.49 259.15 192 ;
      END
   END u2_L10_5_

   PIN u2_L1_23_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 78.85 191.49 78.95 192 ;
      END
   END u2_L1_23_

   PIN u2_L1_28_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 224.85 191.49 224.95 192 ;
      END
   END u2_L1_28_

   PIN u2_L1_9_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 82.95 0.51 83.05 ;
      END
   END u2_L1_9_

   PIN u2_L1_reg_14__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 93.45 191.49 93.55 192 ;
      END
   END u2_L1_reg_14__Q

   PIN u2_L2_18_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.05 191.49 140.15 192 ;
      END
   END u2_L2_18_

   PIN u2_R0_23_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 89.05 191.49 89.15 192 ;
      END
   END u2_R0_23_

   PIN u2_R0_25_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.25 191.49 113.35 192 ;
      END
   END u2_R0_25_

   PIN u2_R0_26_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 202.65 191.49 202.75 192 ;
      END
   END u2_R0_26_

   PIN u2_R0_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 476.25 191.49 476.35 192 ;
      END
   END u2_R0_5_

   PIN u2_R11_15_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 372.25 191.49 372.35 192 ;
      END
   END u2_R11_15_

   PIN u2_R11_21_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 350.25 191.49 350.35 192 ;
      END
   END u2_R11_21_

   PIN u2_R11_27_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 365.05 191.49 365.15 192 ;
      END
   END u2_R11_27_

   PIN u2_R12_22_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 488.45 191.49 488.55 192 ;
      END
   END u2_R12_22_

   PIN u2_R12_28_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 199.65 191.49 199.75 192 ;
      END
   END u2_R12_28_

   PIN u2_R13_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 164.25 191.49 164.35 192 ;
      END
   END u2_R13_5_

   PIN u2_R1_14_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 163.85 191.49 163.95 192 ;
      END
   END u2_R1_14_

   PIN u2_R1_30_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 169.45 191.49 169.55 192 ;
      END
   END u2_R1_30_

   PIN u2_R2_1_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 223.65 191.49 223.75 192 ;
      END
   END u2_R2_1_

   PIN u2_R2_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.85 191.49 67.95 192 ;
      END
   END u2_R2_3_

   PIN u2_R2_6_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.85 191.49 211.95 192 ;
      END
   END u2_R2_6_

   PIN u2_R2_7_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 370.45 191.49 370.55 192 ;
      END
   END u2_R2_7_

   PIN u2_key_r_2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 187.65 191.49 187.75 192 ;
      END
   END u2_key_r_2_

   PIN u2_key_r_35_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 259.25 191.49 259.35 192 ;
      END
   END u2_key_r_35_

   PIN u2_key_r_55_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 176.85 191.49 176.95 192 ;
      END
   END u2_key_r_55_

   PIN u2_key_r_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 142.25 191.49 142.35 192 ;
      END
   END u2_key_r_5_

   PIN u2_uk_K_r_241
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 224.85 191.49 224.95 192 ;
      END
   END u2_uk_K_r_241

   PIN u2_uk_K_r_270
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.05 191.49 80.15 192 ;
      END
   END u2_uk_K_r_270

   OBS
      LAYER via4 ;
         RECT 0 0 523 192 ;
      LAYER via1 ;
         RECT 0 0 523 192 ;
      LAYER metal5 ;
         RECT 0 0 523 192 ;
      LAYER metal4 ;
         RECT 0 0 523 192 ;
      LAYER metal3 ;
         RECT 0 0 523 192 ;
      LAYER metal2 ;
         RECT 0 0 523 192 ;
      LAYER metal1 ;
         RECT 0 0 523 192 ;
   END
END h2

MACRO h1
   CLASS BLOCK ;
   FOREIGN h1 ;
   ORIGIN 0 0 ;
   SIZE 333.2 BY 188 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN1117_n_85315
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 291.45 187.49 291.55 188 ;
      END
   END FE_OFN1117_n_85315

   PIN FE_OFN1131_n_83717
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 144.75 333.2 144.85 ;
      END
   END FE_OFN1131_n_83717

   PIN FE_OFN1447_n_87131
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 308.05 187.49 308.15 188 ;
      END
   END FE_OFN1447_n_87131

   PIN FE_OFN171_n_88228
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.85 187.49 255.95 188 ;
      END
   END FE_OFN171_n_88228

   PIN FE_OFN177_n_87818
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.05 187.49 271.15 188 ;
      END
   END FE_OFN177_n_87818

   PIN FE_OFN183_n_87238
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.85 187.49 234.95 188 ;
      END
   END FE_OFN183_n_87238

   PIN FE_OFN2079_n_83196
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 315.45 187.49 315.55 188 ;
      END
   END FE_OFN2079_n_83196

   PIN FE_OFN2128_n_87090
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 256.25 187.49 256.35 188 ;
      END
   END FE_OFN2128_n_87090

   PIN FE_OFN2671_n_16014
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 144.95 333.2 145.05 ;
      END
   END FE_OFN2671_n_16014

   PIN FE_OFN2969_n_15130
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 315.25 187.49 315.35 188 ;
      END
   END FE_OFN2969_n_15130

   PIN FE_OFN4075_n_84990
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.25 187.49 320.35 188 ;
      END
   END FE_OFN4075_n_84990

   PIN g209359_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 196.85 187.49 196.95 188 ;
      END
   END g209359_p

   PIN g210571_p1
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 256.05 187.49 256.15 188 ;
      END
   END g210571_p1

   PIN g210641_p2
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.45 187.49 292.55 188 ;
      END
   END g210641_p2

   PIN g210835_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 269.65 187.49 269.75 188 ;
      END
   END g210835_sb

   PIN g210889_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 94.95 333.2 95.05 ;
      END
   END g210889_p

   PIN g211048_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 97.15 333.2 97.25 ;
      END
   END g211048_p

   PIN g211616_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 157.75 333.2 157.85 ;
      END
   END g211616_p

   PIN g211975_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 256.25 187.49 256.35 188 ;
      END
   END g211975_db

   PIN g212677_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 298.25 187.49 298.35 188 ;
      END
   END g212677_p

   PIN g213393_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 306.05 187.49 306.15 188 ;
      END
   END g213393_p

   PIN g213779_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.65 187.49 319.75 188 ;
      END
   END g213779_p

   PIN g214217_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 318.05 187.49 318.15 188 ;
      END
   END g214217_db

   PIN g214217_sb
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.45 187.49 321.55 188 ;
      END
   END g214217_sb

   PIN g214307_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 147.35 333.2 147.45 ;
      END
   END g214307_p

   PIN g214357_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.05 187.49 281.15 188 ;
      END
   END g214357_da

   PIN g215900_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 127.55 333.2 127.65 ;
      END
   END g215900_p

   PIN g305635_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 54.85 187.49 54.95 188 ;
      END
   END g305635_da

   PIN g305680_da
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.05 187.49 113.15 188 ;
      END
   END g305680_da

   PIN g305680_db
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.25 187.49 113.35 188 ;
      END
   END g305680_db

   PIN key_b_r_3__184
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 38.65 187.49 38.75 188 ;
      END
   END key_b_r_3__184

   PIN key_c_r_11__1306
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 97.65 187.49 97.75 188 ;
      END
   END key_c_r_11__1306

   PIN key_c_r_19__1727
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 185.45 187.49 185.55 188 ;
      END
   END key_c_r_19__1727

   PIN key_c_r_23__2371
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.65 187.49 124.75 188 ;
      END
   END key_c_r_23__2371

   PIN key_c_r_28__2019
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.45 187.49 128.55 188 ;
      END
   END key_c_r_28__2019

   PIN key_c_r_29__2042
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.65 0 320.75 0.51 ;
      END
   END key_c_r_29__2042

   PIN key_c_r_30__2096
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 172.05 187.49 172.15 188 ;
      END
   END key_c_r_30__2096

   PIN key_c_r_31__2167
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 289.25 187.49 289.35 188 ;
      END
   END key_c_r_31__2167

   PIN key_c_r_32__2208
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 11.95 333.2 12.05 ;
      END
   END key_c_r_32__2208

   PIN key_c_r_32__2234
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 291.65 187.49 291.75 188 ;
      END
   END key_c_r_32__2234

   PIN key_c_r_33__17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 258.25 187.49 258.35 188 ;
      END
   END key_c_r_33__17_

   PIN key_c_r_33__29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 273.45 187.49 273.55 188 ;
      END
   END key_c_r_33__29_

   PIN key_c_r_33__41_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 168.95 333.2 169.05 ;
      END
   END key_c_r_33__41_

   PIN key_c_r_5__2758
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 37.65 187.49 37.75 188 ;
      END
   END key_c_r_5__2758

   PIN key_c_r_8__1129
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 31.25 187.49 31.35 188 ;
      END
   END key_c_r_8__1129

   PIN n_117130
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.05 0 257.15 0.51 ;
      END
   END n_117130

   PIN n_117135
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 269.05 0 269.15 0.51 ;
      END
   END n_117135

   PIN n_126115
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 106.75 333.2 106.85 ;
      END
   END n_126115

   PIN n_15020
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 182.15 333.2 182.25 ;
      END
   END n_15020

   PIN n_15309
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 171.95 333.2 172.05 ;
      END
   END n_15309

   PIN n_15373
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.45 187.49 319.55 188 ;
      END
   END n_15373

   PIN n_15376
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 157.95 333.2 158.05 ;
      END
   END n_15376

   PIN n_15814
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.85 187.49 321.95 188 ;
      END
   END n_15814

   PIN n_16235
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 145.15 333.2 145.25 ;
      END
   END n_16235

   PIN n_16236
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 172.15 333.2 172.25 ;
      END
   END n_16236

   PIN n_599
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 135.05 187.49 135.15 188 ;
      END
   END n_599

   PIN n_636
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 48.85 187.49 48.95 188 ;
      END
   END n_636

   PIN n_643
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 89.05 187.49 89.15 188 ;
      END
   END n_643

   PIN n_82873
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 112.35 333.2 112.45 ;
      END
   END n_82873

   PIN n_82885
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 131.95 333.2 132.05 ;
      END
   END n_82885

   PIN n_82988
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 305.85 187.49 305.95 188 ;
      END
   END n_82988

   PIN n_83094
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 120.55 333.2 120.65 ;
      END
   END n_83094

   PIN n_83137
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 147.35 333.2 147.45 ;
      END
   END n_83137

   PIN n_83203
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 269.05 187.49 269.15 188 ;
      END
   END n_83203

   PIN n_83256
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 121.35 333.2 121.45 ;
      END
   END n_83256

   PIN n_83274
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 141.35 333.2 141.45 ;
      END
   END n_83274

   PIN n_83283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 122.75 333.2 122.85 ;
      END
   END n_83283

   PIN n_83296
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 121.55 333.2 121.65 ;
      END
   END n_83296

   PIN n_83307
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 36.15 333.2 36.25 ;
      END
   END n_83307

   PIN n_83371
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 108.15 333.2 108.25 ;
      END
   END n_83371

   PIN n_83404
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 116.55 333.2 116.65 ;
      END
   END n_83404

   PIN n_83450
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 119.75 333.2 119.85 ;
      END
   END n_83450

   PIN n_83520
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 119.15 333.2 119.25 ;
      END
   END n_83520

   PIN n_83598
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 122.15 333.2 122.25 ;
      END
   END n_83598

   PIN n_83639
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 156.35 333.2 156.45 ;
      END
   END n_83639

   PIN n_83663
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 120.95 333.2 121.05 ;
      END
   END n_83663

   PIN n_83674
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 24.75 333.2 24.85 ;
      END
   END n_83674

   PIN n_83733
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 130.15 333.2 130.25 ;
      END
   END n_83733

   PIN n_83783
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 124.55 333.2 124.65 ;
      END
   END n_83783

   PIN n_83805
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.65 0 320.75 0.51 ;
      END
   END n_83805

   PIN n_83907
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 141.15 333.2 141.25 ;
      END
   END n_83907

   PIN n_83923
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 23.95 333.2 24.05 ;
      END
   END n_83923

   PIN n_83974
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 118.95 333.2 119.05 ;
      END
   END n_83974

   PIN n_84019
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 145.75 333.2 145.85 ;
      END
   END n_84019

   PIN n_84035
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 120.75 333.2 120.85 ;
      END
   END n_84035

   PIN n_84063
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 130.35 333.2 130.45 ;
      END
   END n_84063

   PIN n_84124
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 121.75 333.2 121.85 ;
      END
   END n_84124

   PIN n_84128
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 125.55 333.2 125.65 ;
      END
   END n_84128

   PIN n_84129
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 125.75 333.2 125.85 ;
      END
   END n_84129

   PIN n_84154
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 107.75 333.2 107.85 ;
      END
   END n_84154

   PIN n_84252
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 123.55 333.2 123.65 ;
      END
   END n_84252

   PIN n_84301
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 107.95 333.2 108.05 ;
      END
   END n_84301

   PIN n_84317
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 107.35 333.2 107.45 ;
      END
   END n_84317

   PIN n_84327
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 121.95 333.2 122.05 ;
      END
   END n_84327

   PIN n_84402
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 121.55 333.2 121.65 ;
      END
   END n_84402

   PIN n_84435
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 140.75 333.2 140.85 ;
      END
   END n_84435

   PIN n_84440
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 127.75 333.2 127.85 ;
      END
   END n_84440

   PIN n_84544
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 112.15 333.2 112.25 ;
      END
   END n_84544

   PIN n_84557
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 124.75 333.2 124.85 ;
      END
   END n_84557

   PIN n_84593
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 132.95 333.2 133.05 ;
      END
   END n_84593

   PIN n_84597
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 130.75 333.2 130.85 ;
      END
   END n_84597

   PIN n_84610
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 107.55 333.2 107.65 ;
      END
   END n_84610

   PIN n_84652
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.45 0 320.55 0.51 ;
      END
   END n_84652

   PIN n_84873
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 138.95 333.2 139.05 ;
      END
   END n_84873

   PIN n_84915
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 151.75 333.2 151.85 ;
      END
   END n_84915

   PIN n_84933
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 141.95 333.2 142.05 ;
      END
   END n_84933

   PIN n_84971
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 139.15 333.2 139.25 ;
      END
   END n_84971

   PIN n_84986
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 156.55 333.2 156.65 ;
      END
   END n_84986

   PIN n_84988
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 139.35 333.2 139.45 ;
      END
   END n_84988

   PIN n_84998
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 291.85 187.49 291.95 188 ;
      END
   END n_84998

   PIN n_84999
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 141.55 333.2 141.65 ;
      END
   END n_84999

   PIN n_85002
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 168.15 333.2 168.25 ;
      END
   END n_85002

   PIN n_85013
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 148.95 333.2 149.05 ;
      END
   END n_85013

   PIN n_85031
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 153.15 333.2 153.25 ;
      END
   END n_85031

   PIN n_85033
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 137.75 333.2 137.85 ;
      END
   END n_85033

   PIN n_85037
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 144.95 333.2 145.05 ;
      END
   END n_85037

   PIN n_85044
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 116.75 333.2 116.85 ;
      END
   END n_85044

   PIN n_85059
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.85 187.49 220.95 188 ;
      END
   END n_85059

   PIN n_85086
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.65 187.49 320.75 188 ;
      END
   END n_85086

   PIN n_85103
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 294.45 187.49 294.55 188 ;
      END
   END n_85103

   PIN n_85147
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 305.65 187.49 305.75 188 ;
      END
   END n_85147

   PIN n_85176
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.05 187.49 282.15 188 ;
      END
   END n_85176

   PIN n_85187
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 145.15 333.2 145.25 ;
      END
   END n_85187

   PIN n_85208
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 151.95 333.2 152.05 ;
      END
   END n_85208

   PIN n_85249
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 292.05 187.49 292.15 188 ;
      END
   END n_85249

   PIN n_85270
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 306.85 187.49 306.95 188 ;
      END
   END n_85270

   PIN n_85275
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 156.75 333.2 156.85 ;
      END
   END n_85275

   PIN n_85344
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.945 155.3 333.2 155.5 ;
      END
   END n_85344

   PIN n_85378
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.25 187.49 258.35 188 ;
      END
   END n_85378

   PIN n_85405
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 280.65 187.49 280.75 188 ;
      END
   END n_85405

   PIN n_85406
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.65 187.49 294.75 188 ;
      END
   END n_85406

   PIN n_85475
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 279.65 187.49 279.75 188 ;
      END
   END n_85475

   PIN n_85559
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 170.35 333.2 170.45 ;
      END
   END n_85559

   PIN n_85684
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 270.2 187.745 270.4 188 ;
      END
   END n_85684

   PIN n_85696
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.25 187.49 282.35 188 ;
      END
   END n_85696

   PIN n_85699
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 267.85 187.49 267.95 188 ;
      END
   END n_85699

   PIN n_85700
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 269.25 187.49 269.35 188 ;
      END
   END n_85700

   PIN n_85722
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 155.95 333.2 156.05 ;
      END
   END n_85722

   PIN n_85818
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.85 187.49 283.95 188 ;
      END
   END n_85818

   PIN n_85821
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.25 187.49 281.35 188 ;
      END
   END n_85821

   PIN n_85842
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.85 187.49 270.95 188 ;
      END
   END n_85842

   PIN n_85870
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 154.95 333.2 155.05 ;
      END
   END n_85870

   PIN n_85877
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 168.55 333.2 168.65 ;
      END
   END n_85877

   PIN n_85878
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 168.75 333.2 168.85 ;
      END
   END n_85878

   PIN n_85879
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 167.95 333.2 168.05 ;
      END
   END n_85879

   PIN n_85946
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 225.05 187.49 225.15 188 ;
      END
   END n_85946

   PIN n_85967
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 154.75 333.2 154.85 ;
      END
   END n_85967

   PIN n_85970
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 292.25 187.49 292.35 188 ;
      END
   END n_85970

   PIN n_85991
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 156.35 333.2 156.45 ;
      END
   END n_85991

   PIN n_86002
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 182.35 333.2 182.45 ;
      END
   END n_86002

   PIN n_86110
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.65 187.49 271.75 188 ;
      END
   END n_86110

   PIN n_86119
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 269.05 187.49 269.15 188 ;
      END
   END n_86119

   PIN n_86129
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 154.35 333.2 154.45 ;
      END
   END n_86129

   PIN n_86135
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.45 187.49 283.55 188 ;
      END
   END n_86135

   PIN n_86142
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 181.35 333.2 181.45 ;
      END
   END n_86142

   PIN n_86146
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 182.55 333.2 182.65 ;
      END
   END n_86146

   PIN n_86151
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 141.95 333.2 142.05 ;
      END
   END n_86151

   PIN n_86152
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 292.45 187.49 292.55 188 ;
      END
   END n_86152

   PIN n_86238
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 269.25 187.49 269.35 188 ;
      END
   END n_86238

   PIN n_86246
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.25 187.49 271.35 188 ;
      END
   END n_86246

   PIN n_86249
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 154.15 333.2 154.25 ;
      END
   END n_86249

   PIN n_86258
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 170.55 333.2 170.65 ;
      END
   END n_86258

   PIN n_86296
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 168.95 333.2 169.05 ;
      END
   END n_86296

   PIN n_86305
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 172.35 333.2 172.45 ;
      END
   END n_86305

   PIN n_86355
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 109.95 333.2 110.05 ;
      END
   END n_86355

   PIN n_86362
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.65 187.49 292.75 188 ;
      END
   END n_86362

   PIN n_86364
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 305.05 187.49 305.15 188 ;
      END
   END n_86364

   PIN n_86365
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 257.8 187.745 258 188 ;
      END
   END n_86365

   PIN n_86383
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 168.75 333.2 168.85 ;
      END
   END n_86383

   PIN n_86431
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 182.75 333.2 182.85 ;
      END
   END n_86431

   PIN n_86433
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 103.95 333.2 104.05 ;
      END
   END n_86433

   PIN n_86440
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.45 187.49 281.55 188 ;
      END
   END n_86440

   PIN n_86479
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.25 187.49 292.35 188 ;
      END
   END n_86479

   PIN n_86494
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 279.85 187.49 279.95 188 ;
      END
   END n_86494

   PIN n_86540
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 294.65 187.49 294.75 188 ;
      END
   END n_86540

   PIN n_86551
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 172.55 333.2 172.65 ;
      END
   END n_86551

   PIN n_86592
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 269.45 187.49 269.55 188 ;
      END
   END n_86592

   PIN n_86600
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 256.45 187.49 256.55 188 ;
      END
   END n_86600

   PIN n_86621
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.05 187.49 197.15 188 ;
      END
   END n_86621

   PIN n_86643
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 300.05 187.49 300.15 188 ;
      END
   END n_86643

   PIN n_86645
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 168.15 333.2 168.25 ;
      END
   END n_86645

   PIN n_86646
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 298.05 187.49 298.15 188 ;
      END
   END n_86646

   PIN n_86674
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.25 187.49 197.35 188 ;
      END
   END n_86674

   PIN n_86688
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 305.25 187.49 305.35 188 ;
      END
   END n_86688

   PIN n_86724
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 300.85 187.49 300.95 188 ;
      END
   END n_86724

   PIN n_86745
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 197.05 187.49 197.15 188 ;
      END
   END n_86745

   PIN n_86793
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 133.15 333.2 133.25 ;
      END
   END n_86793

   PIN n_86805
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 293.45 187.49 293.55 188 ;
      END
   END n_86805

   PIN n_86808
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 107.15 333.2 107.25 ;
      END
   END n_86808

   PIN n_86828
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 156.95 333.2 157.05 ;
      END
   END n_86828

   PIN n_86842
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 153.35 333.2 153.45 ;
      END
   END n_86842

   PIN n_86858
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 143.15 333.2 143.25 ;
      END
   END n_86858

   PIN n_87007
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 156.75 333.2 156.85 ;
      END
   END n_87007

   PIN n_87056
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 149.35 333.2 149.45 ;
      END
   END n_87056

   PIN n_87144
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 234.45 187.49 234.55 188 ;
      END
   END n_87144

   PIN n_87202
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 295.85 187.49 295.95 188 ;
      END
   END n_87202

   PIN n_87212
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 282.45 187.49 282.55 188 ;
      END
   END n_87212

   PIN n_87219
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.945 71.7 333.2 71.9 ;
      END
   END n_87219

   PIN n_87221
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 184.85 187.49 184.95 188 ;
      END
   END n_87221

   PIN n_87239
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 245.85 187.49 245.95 188 ;
      END
   END n_87239

   PIN n_87240
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 256.45 187.49 256.55 188 ;
      END
   END n_87240

   PIN n_87294
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.05 187.49 233.15 188 ;
      END
   END n_87294

   PIN n_87311
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 246.6 187.745 246.8 188 ;
      END
   END n_87311

   PIN n_87321
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 99.35 333.2 99.45 ;
      END
   END n_87321

   PIN n_87330
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 148.85 187.49 148.95 188 ;
      END
   END n_87330

   PIN n_87336
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 271.45 187.49 271.55 188 ;
      END
   END n_87336

   PIN n_87368
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.65 187.49 258.75 188 ;
      END
   END n_87368

   PIN n_87394
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 295.05 187.49 295.15 188 ;
      END
   END n_87394

   PIN n_87399
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.25 187.49 233.35 188 ;
      END
   END n_87399

   PIN n_87412
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.65 187.49 234.75 188 ;
      END
   END n_87412

   PIN n_87421
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.65 187.49 245.75 188 ;
      END
   END n_87421

   PIN n_87424
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 69.15 333.2 69.25 ;
      END
   END n_87424

   PIN n_87472
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.945 148.1 333.2 148.3 ;
      END
   END n_87472

   PIN n_87486
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 69.35 333.2 69.45 ;
      END
   END n_87486

   PIN n_87498
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 246.25 187.49 246.35 188 ;
      END
   END n_87498

   PIN n_87530
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 234.65 187.49 234.75 188 ;
      END
   END n_87530

   PIN n_87556
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 246.05 187.49 246.15 188 ;
      END
   END n_87556

   PIN n_87572
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 232.25 187.49 232.35 188 ;
      END
   END n_87572

   PIN n_87580
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 294.85 187.49 294.95 188 ;
      END
   END n_87580

   PIN n_87586
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 225.25 187.49 225.35 188 ;
      END
   END n_87586

   PIN n_87593
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 94.35 333.2 94.45 ;
      END
   END n_87593

   PIN n_87600
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 256.65 187.49 256.75 188 ;
      END
   END n_87600

   PIN n_87616
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 269.45 187.49 269.55 188 ;
      END
   END n_87616

   PIN n_87642
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 69.55 333.2 69.65 ;
      END
   END n_87642

   PIN n_87644
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 257.05 187.49 257.15 188 ;
      END
   END n_87644

   PIN n_87648
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 124.85 187.49 124.95 188 ;
      END
   END n_87648

   PIN n_87657
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 94.55 333.2 94.65 ;
      END
   END n_87657

   PIN n_87697
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 295.4 187.745 295.6 188 ;
      END
   END n_87697

   PIN n_87745
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285.65 187.49 285.75 188 ;
      END
   END n_87745

   PIN n_87752
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.65 187.49 281.75 188 ;
      END
   END n_87752

   PIN n_87753
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 269.85 187.49 269.95 188 ;
      END
   END n_87753

   PIN n_87757
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.05 187.49 307.15 188 ;
      END
   END n_87757

   PIN n_87789
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 172.85 187.49 172.95 188 ;
      END
   END n_87789

   PIN n_87794
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.65 187.49 293.75 188 ;
      END
   END n_87794

   PIN n_87812
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.45 187.49 233.55 188 ;
      END
   END n_87812

   PIN n_87816
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 306.45 187.49 306.55 188 ;
      END
   END n_87816

   PIN n_87818
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 85.15 333.2 85.25 ;
      END
   END n_87818

   PIN n_87821
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.25 187.49 221.35 188 ;
      END
   END n_87821

   PIN n_87839
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.05 187.49 221.15 188 ;
      END
   END n_87839

   PIN n_87875
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.45 187.49 258.55 188 ;
      END
   END n_87875

   PIN n_87932
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 256.85 187.49 256.95 188 ;
      END
   END n_87932

   PIN n_87934
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.945 130.7 333.2 130.9 ;
      END
   END n_87934

   PIN n_87935
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 209.25 187.49 209.35 188 ;
      END
   END n_87935

   PIN n_87944
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 225.45 187.49 225.55 188 ;
      END
   END n_87944

   PIN n_87945
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 197.45 187.49 197.55 188 ;
      END
   END n_87945

   PIN n_87951
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.45 187.49 257.55 188 ;
      END
   END n_87951

   PIN n_88028
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 268.05 187.49 268.15 188 ;
      END
   END n_88028

   PIN n_88056
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 317.45 187.49 317.55 188 ;
      END
   END n_88056

   PIN n_88065
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285.25 187.49 285.35 188 ;
      END
   END n_88065

   PIN n_88067
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 322.05 187.49 322.15 188 ;
      END
   END n_88067

   PIN n_88085
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 269.65 187.49 269.75 188 ;
      END
   END n_88085

   PIN n_88092
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 281.85 187.49 281.95 188 ;
      END
   END n_88092

   PIN n_88094
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 293.65 187.49 293.75 188 ;
      END
   END n_88094

   PIN n_88111
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 246.65 187.49 246.75 188 ;
      END
   END n_88111

   PIN n_88115
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.25 187.49 307.35 188 ;
      END
   END n_88115

   PIN n_88121
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 173.05 187.49 173.15 188 ;
      END
   END n_88121

   PIN n_88124
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.85 187.49 293.95 188 ;
      END
   END n_88124

   PIN n_88191
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 142.75 333.2 142.85 ;
      END
   END n_88191

   PIN n_88200
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 268.25 187.49 268.35 188 ;
      END
   END n_88200

   PIN n_88216
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 295.05 187.49 295.15 188 ;
      END
   END n_88216

   PIN n_88257
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 88.95 333.2 89.05 ;
      END
   END n_88257

   PIN n_88341
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 318.25 187.49 318.35 188 ;
      END
   END n_88341

   PIN n_88342
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 99.15 333.2 99.25 ;
      END
   END n_88342

   PIN n_88348
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.05 187.49 294.15 188 ;
      END
   END n_88348

   PIN n_88351
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.85 187.49 258.95 188 ;
      END
   END n_88351

   PIN n_88352
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 269.85 187.49 269.95 188 ;
      END
   END n_88352

   PIN n_88358
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 280.05 187.49 280.15 188 ;
      END
   END n_88358

   PIN n_88359
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 97.35 333.2 97.45 ;
      END
   END n_88359

   PIN n_88383
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 268.45 187.49 268.55 188 ;
      END
   END n_88383

   PIN n_88433
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 292.65 187.49 292.75 188 ;
      END
   END n_88433

   PIN n_88466
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.65 187.49 257.75 188 ;
      END
   END n_88466

   PIN n_88505
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 256.65 187.49 256.75 188 ;
      END
   END n_88505

   PIN n_88508
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 256.85 187.49 256.95 188 ;
      END
   END n_88508

   PIN n_88519
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 280.25 187.49 280.35 188 ;
      END
   END n_88519

   PIN n_88570
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.05 187.49 245.15 188 ;
      END
   END n_88570

   PIN n_88591
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.05 187.49 257.15 188 ;
      END
   END n_88591

   PIN n_88603
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 101.15 333.2 101.25 ;
      END
   END n_88603

   PIN n_88633
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.85 187.49 319.95 188 ;
      END
   END n_88633

   PIN n_88640
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 232.45 187.49 232.55 188 ;
      END
   END n_88640

   PIN n_88657
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.85 187.49 294.95 188 ;
      END
   END n_88657

   PIN n_88669
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 257.25 187.49 257.35 188 ;
      END
   END n_88669

   PIN n_88670
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.25 187.49 319.35 188 ;
      END
   END n_88670

   PIN n_88681
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 292.85 187.49 292.95 188 ;
      END
   END n_88681

   PIN n_88726
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 135.35 333.2 135.45 ;
      END
   END n_88726

   PIN n_88770
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 306.65 187.49 306.75 188 ;
      END
   END n_88770

   PIN n_88771
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 315.05 187.49 315.15 188 ;
      END
   END n_88771

   PIN n_88781
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 233.65 187.49 233.75 188 ;
      END
   END n_88781

   PIN n_88782
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 232.65 187.49 232.75 188 ;
      END
   END n_88782

   PIN n_88793
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 132.95 333.2 133.05 ;
      END
   END n_88793

   PIN n_88815
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 59.95 333.2 60.05 ;
      END
   END n_88815

   PIN n_88816
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 306.25 187.49 306.35 188 ;
      END
   END n_88816

   PIN n_88842
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 308.25 187.49 308.35 188 ;
      END
   END n_88842

   PIN n_88874
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 71.35 333.2 71.45 ;
      END
   END n_88874

   PIN n_88877
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 305.45 187.49 305.55 188 ;
      END
   END n_88877

   PIN n_88897
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 127.95 333.2 128.05 ;
      END
   END n_88897

   PIN n_89163
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 313.25 187.49 313.35 188 ;
      END
   END n_89163

   PIN n_89299
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 293.85 187.49 293.95 188 ;
      END
   END n_89299

   PIN n_89430
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 158.15 333.2 158.25 ;
      END
   END n_89430

   PIN n_89487
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 304.85 187.49 304.95 188 ;
      END
   END n_89487

   PIN n_89527
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.45 187.49 221.55 188 ;
      END
   END n_89527

   PIN n_89607
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 145.95 333.2 146.05 ;
      END
   END n_89607

   PIN n_89612
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 310.05 187.49 310.15 188 ;
      END
   END n_89612

   PIN n_89671
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 311.05 187.49 311.15 188 ;
      END
   END n_89671

   PIN n_89743
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 138.75 333.2 138.85 ;
      END
   END n_89743

   PIN n_89790
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 314.65 187.49 314.75 188 ;
      END
   END n_89790

   PIN n_89829
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.45 187.49 308.55 188 ;
      END
   END n_89829

   PIN n_89924
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 182.95 333.2 183.05 ;
      END
   END n_89924

   PIN n_89926
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 168.35 333.2 168.45 ;
      END
   END n_89926

   PIN n_89927
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 268.65 187.49 268.75 188 ;
      END
   END n_89927

   PIN n_89999
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 317.45 187.49 317.55 188 ;
      END
   END n_89999

   PIN n_90006
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 144.55 333.2 144.65 ;
      END
   END n_90006

   PIN n_90059
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.85 187.49 306.95 188 ;
      END
   END n_90059

   PIN n_90215
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 294.05 187.49 294.15 188 ;
      END
   END n_90215

   PIN n_90279
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 309.85 187.49 309.95 188 ;
      END
   END n_90279

   PIN n_90333
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 309.45 187.49 309.55 188 ;
      END
   END n_90333

   PIN n_90412
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 309.45 187.49 309.55 188 ;
      END
   END n_90412

   PIN n_90417
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 317.65 187.49 317.75 188 ;
      END
   END n_90417

   PIN n_90560
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 209.45 187.49 209.55 188 ;
      END
   END n_90560

   PIN n_90687
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 315.65 187.49 315.75 188 ;
      END
   END n_90687

   PIN n_90693
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 183.15 333.2 183.25 ;
      END
   END n_90693

   PIN n_90818
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 136.75 333.2 136.85 ;
      END
   END n_90818

   PIN n_90859
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 139.55 333.2 139.65 ;
      END
   END n_90859

   PIN u1_key_r_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 236.25 187.49 236.35 188 ;
      END
   END u1_key_r_2_

   PIN u1_key_r_30_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285.85 187.49 285.95 188 ;
      END
   END u1_key_r_30_

   PIN u1_key_r_55_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 250.05 187.49 250.15 188 ;
      END
   END u1_key_r_55_

   PIN u2_L2_17_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 139.75 333.2 139.85 ;
      END
   END u2_L2_17_

   PIN u2_L3_18_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.65 187.49 221.75 188 ;
      END
   END u2_L3_18_

   PIN u2_L3_reg_14__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.05 187.49 319.15 188 ;
      END
   END u2_L3_reg_14__Q

   PIN u2_L4_18_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 145.55 333.2 145.65 ;
      END
   END u2_L4_18_

   PIN u2_L4_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 136.55 333.2 136.65 ;
      END
   END u2_L4_28_

   PIN u2_L4_32_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.65 187.49 233.75 188 ;
      END
   END u2_L4_32_

   PIN u2_L4_8_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 232.85 187.49 232.95 188 ;
      END
   END u2_L4_8_

   PIN u2_L5_14_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 139.95 333.2 140.05 ;
      END
   END u2_L5_14_

   PIN u2_L5_30_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 318.85 187.49 318.95 188 ;
      END
   END u2_L5_30_

   PIN u2_L5_reg_12__Q
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 140.15 333.2 140.25 ;
      END
   END u2_L5_reg_12__Q

   PIN u2_R3_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.05 0 293.15 0.51 ;
      END
   END u2_R3_1_

   PIN u2_R3_2_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 319.45 187.49 319.55 188 ;
      END
   END u2_R3_2_

   PIN u2_R3_7_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 128.15 333.2 128.25 ;
      END
   END u2_R3_7_

   PIN u2_R4_13_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 257.45 187.49 257.55 188 ;
      END
   END u2_R4_13_

   PIN u2_R4_22_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 156.15 333.2 156.25 ;
      END
   END u2_R4_22_

   PIN u2_R4_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 183.35 333.2 183.45 ;
      END
   END u2_R4_23_

   PIN u2_R4_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.05 187.49 270.15 188 ;
      END
   END u2_R4_28_

   PIN u2_R4_29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 145.35 333.2 145.45 ;
      END
   END u2_R4_29_

   PIN u2_R4_3_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 293.05 187.49 293.15 188 ;
      END
   END u2_R4_3_

   PIN u2_R5_12_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 119.35 333.2 119.45 ;
      END
   END u2_R5_12_

   PIN u2_R5_29_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 116.95 333.2 117.05 ;
      END
   END u2_R5_29_

   PIN u2_R5_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 60.15 333.2 60.25 ;
      END
   END u2_R5_4_

   PIN u2_key_r_21_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 222.05 187.49 222.15 188 ;
      END
   END u2_key_r_21_

   PIN u2_uk_K_r_530
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 138.55 333.2 138.65 ;
      END
   END u2_uk_K_r_530

   PIN FE_OFN1065_n_116
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 291 187.745 291.2 188 ;
      END
   END FE_OFN1065_n_116

   PIN FE_OFN1130_n_82876
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 133.15 333.2 133.25 ;
      END
   END FE_OFN1130_n_82876

   PIN FE_OFN1354_n_88664
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 154.35 333.2 154.45 ;
      END
   END FE_OFN1354_n_88664

   PIN FE_OFN1476_n_15154
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 129.95 333.2 130.05 ;
      END
   END FE_OFN1476_n_15154

   PIN FE_OFN1597_n_16688
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 115.95 333.2 116.05 ;
      END
   END FE_OFN1597_n_16688

   PIN FE_OFN176_n_87818
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 84.95 333.2 85.05 ;
      END
   END FE_OFN176_n_87818

   PIN FE_OFN1837_n_16002
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 130.95 333.2 131.05 ;
      END
   END FE_OFN1837_n_16002

   PIN FE_OFN1909_n_85016
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 147.15 333.2 147.25 ;
      END
   END FE_OFN1909_n_85016

   PIN FE_OFN2000_n_84960
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 128.75 333.2 128.85 ;
      END
   END FE_OFN2000_n_84960

   PIN FE_OFN2127_n_87090
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 232.05 187.49 232.15 188 ;
      END
   END FE_OFN2127_n_87090

   PIN FE_OFN2410_n_82958
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 180.15 333.2 180.25 ;
      END
   END FE_OFN2410_n_82958

   PIN FE_OFN2514_n_82929
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.945 124.1 333.2 124.3 ;
      END
   END FE_OFN2514_n_82929

   PIN FE_OFN2809_n_16012
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 181.15 333.2 181.25 ;
      END
   END FE_OFN2809_n_16012

   PIN FE_OFN2888_n_16011
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 314.25 187.49 314.35 188 ;
      END
   END FE_OFN2888_n_16011

   PIN FE_OFN3132_n_16013
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 134.95 333.2 135.05 ;
      END
   END FE_OFN3132_n_16013

   PIN FE_OFN3225_n_15131
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 146.95 333.2 147.05 ;
      END
   END FE_OFN3225_n_15131

   PIN FE_OFN3320_n_500
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 50 187.745 50.2 188 ;
      END
   END FE_OFN3320_n_500

   PIN FE_OFN3436_n_89910
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 310.65 187.49 310.75 188 ;
      END
   END FE_OFN3436_n_89910

   PIN FE_OFN3698_n_16007
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.45 187.49 307.55 188 ;
      END
   END FE_OFN3698_n_16007

   PIN FE_OFN4024_n_85019
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 133.95 333.2 134.05 ;
      END
   END FE_OFN4024_n_85019

   PIN FE_OFN4400_decrypt
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.945 155.1 333.2 155.3 ;
      END
   END FE_OFN4400_decrypt

   PIN FE_OFN4722_n_500
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 233.2 187.745 233.4 188 ;
      END
   END FE_OFN4722_n_500

   PIN FE_OFN4816_n_16014
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 171.75 333.2 171.85 ;
      END
   END FE_OFN4816_n_16014

   PIN FE_OFN872_n_84986
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 156.95 333.2 157.05 ;
      END
   END FE_OFN872_n_84986

   PIN g210626_p1
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.45 187.49 232.55 188 ;
      END
   END g210626_p1

   PIN g210918_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.45 187.49 318.55 188 ;
      END
   END g210918_p

   PIN g211000_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 209.05 187.49 209.15 188 ;
      END
   END g211000_p

   PIN g211245_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 149.15 333.2 149.25 ;
      END
   END g211245_p

   PIN g211261_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 74.95 333.2 75.05 ;
      END
   END g211261_p

   PIN g211472_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 256.05 187.49 256.15 188 ;
      END
   END g211472_p

   PIN g211617_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 220.65 187.49 220.75 188 ;
      END
   END g211617_p

   PIN g211748_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.05 187.49 292.15 188 ;
      END
   END g211748_p

   PIN g212987_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 268.85 187.49 268.95 188 ;
      END
   END g212987_p

   PIN g214406_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 309.05 187.49 309.15 188 ;
      END
   END g214406_db

   PIN g214423_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 137.55 333.2 137.65 ;
      END
   END g214423_db

   PIN g214423_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 135.15 333.2 135.25 ;
      END
   END g214423_sb

   PIN g216122_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 144.55 333.2 144.65 ;
      END
   END g216122_sb

   PIN g216695_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 315.05 187.49 315.15 188 ;
      END
   END g216695_sb

   PIN g286480_p
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 171.55 333.2 171.65 ;
      END
   END g286480_p

   PIN g305627_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.25 187.49 55.35 188 ;
      END
   END g305627_sb

   PIN g305634_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 65.05 187.49 65.15 188 ;
      END
   END g305634_da

   PIN g305634_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.05 187.49 52.15 188 ;
      END
   END g305634_db

   PIN g305715_da
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 49.05 187.49 49.15 188 ;
      END
   END g305715_da

   PIN g321810_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.65 187.49 255.75 188 ;
      END
   END g321810_db

   PIN g321810_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.45 187.49 255.55 188 ;
      END
   END g321810_sb

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.945 132.3 333.2 132.5 ;
      END
   END ispd_clk

   PIN key1_17_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 55.05 187.49 55.15 188 ;
      END
   END key1_17_

   PIN key1_37_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 135.65 187.49 135.75 188 ;
      END
   END key1_37_

   PIN key1_39_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.85 187.49 232.95 188 ;
      END
   END key1_39_

   PIN key2_19_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 132.15 0.51 132.25 ;
      END
   END key2_19_

   PIN key3_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 45.25 187.49 45.35 188 ;
      END
   END key3_11_

   PIN key3_37_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 52.45 187.49 52.55 188 ;
      END
   END key3_37_

   PIN key3_39_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.65 187.49 232.75 188 ;
      END
   END key3_39_

   PIN key_b_r_15__880
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 147.05 187.49 147.15 188 ;
      END
   END key_b_r_15__880

   PIN key_b_r_16__2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.65 187.49 29.75 188 ;
      END
   END key_b_r_16__2_

   PIN key_b_r_16__30_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 40.85 187.49 40.95 188 ;
      END
   END key_b_r_16__30_

   PIN key_c_r_20__1782
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 196.65 187.49 196.75 188 ;
      END
   END key_c_r_20__1782

   PIN key_c_r_21__1822
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.45 187.49 29.55 188 ;
      END
   END key_c_r_21__1822

   PIN key_c_r_27__1931
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 157.45 187.49 157.55 188 ;
      END
   END key_c_r_27__1931

   PIN key_c_r_27__1964
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.85 187.49 112.95 188 ;
      END
   END key_c_r_27__1964

   PIN key_c_r_27__1966
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 112.65 187.49 112.75 188 ;
      END
   END key_c_r_27__1966

   PIN key_c_r_2__2648
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 22.25 187.49 22.35 188 ;
      END
   END key_c_r_2__2648

   PIN key_c_r_30__2098
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.25 187.49 77.35 188 ;
      END
   END key_c_r_30__2098

   PIN key_c_r_31__2162
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 17.05 187.49 17.15 188 ;
      END
   END key_c_r_31__2162

   PIN key_c_r_31__2179
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 77.05 187.49 77.15 188 ;
      END
   END key_c_r_31__2179

   PIN key_c_r_32__2221
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.25 187.49 29.35 188 ;
      END
   END key_c_r_32__2221

   PIN key_c_r_32__2229
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 76.85 187.49 76.95 188 ;
      END
   END key_c_r_32__2229

   PIN key_c_r_5__2791
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 29.05 187.49 29.15 188 ;
      END
   END key_c_r_5__2791

   PIN key_c_r_6__1019
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 17.05 187.49 17.15 188 ;
      END
   END key_c_r_6__1019

   PIN key_c_r_7__1051
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 105.45 187.49 105.55 188 ;
      END
   END key_c_r_7__1051

   PIN key_c_r_9__1177
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 113.45 187.49 113.55 188 ;
      END
   END key_c_r_9__1177

   PIN n_108924
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 268.65 187.49 268.75 188 ;
      END
   END n_108924

   PIN n_108925
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.25 187.49 255.35 188 ;
      END
   END n_108925

   PIN n_118831
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 305.45 187.49 305.55 188 ;
      END
   END n_118831

   PIN n_118867
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 209.05 187.49 209.15 188 ;
      END
   END n_118867

   PIN n_14583
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 181.95 333.2 182.05 ;
      END
   END n_14583

   PIN n_15021
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 137.35 333.2 137.45 ;
      END
   END n_15021

   PIN n_15130
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 144.35 333.2 144.45 ;
      END
   END n_15130

   PIN n_15136
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 316.25 187.49 316.35 188 ;
      END
   END n_15136

   PIN n_15152
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 315.85 187.49 315.95 188 ;
      END
   END n_15152

   PIN n_15372
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 316.45 187.49 316.55 188 ;
      END
   END n_15372

   PIN n_15780
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 171.35 333.2 171.45 ;
      END
   END n_15780

   PIN n_15789
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 181.75 333.2 181.85 ;
      END
   END n_15789

   PIN n_15811
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 317.05 187.49 317.15 188 ;
      END
   END n_15811

   PIN n_15813
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 170.15 333.2 170.25 ;
      END
   END n_15813

   PIN n_15820
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 169.95 333.2 170.05 ;
      END
   END n_15820

   PIN n_15823
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 180.95 333.2 181.05 ;
      END
   END n_15823

   PIN n_15989
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 128.95 333.2 129.05 ;
      END
   END n_15989

   PIN n_16001
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 314.45 187.49 314.55 188 ;
      END
   END n_16001

   PIN n_16005
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 168.55 333.2 168.65 ;
      END
   END n_16005

   PIN n_16006
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 140.35 333.2 140.45 ;
      END
   END n_16006

   PIN n_16008
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 318.65 187.49 318.75 188 ;
      END
   END n_16008

   PIN n_16010
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 180.75 333.2 180.85 ;
      END
   END n_16010

   PIN n_16015
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.85 187.49 291.95 188 ;
      END
   END n_16015

   PIN n_16017
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 135.75 333.2 135.85 ;
      END
   END n_16017

   PIN n_16021
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 169.75 333.2 169.85 ;
      END
   END n_16021

   PIN n_16022
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 140.55 333.2 140.65 ;
      END
   END n_16022

   PIN n_16140
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 180.55 333.2 180.65 ;
      END
   END n_16140

   PIN n_16141
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 317.65 187.49 317.75 188 ;
      END
   END n_16141

   PIN n_16195
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 148.95 333.2 149.05 ;
      END
   END n_16195

   PIN n_16229
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 143.35 333.2 143.45 ;
      END
   END n_16229

   PIN n_16233
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.05 187.49 320.15 188 ;
      END
   END n_16233

   PIN n_16511
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 308.85 187.49 308.95 188 ;
      END
   END n_16511

   PIN n_16677
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 180.35 333.2 180.45 ;
      END
   END n_16677

   PIN n_16679
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 147.75 333.2 147.85 ;
      END
   END n_16679

   PIN n_16680
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.85 187.49 319.95 188 ;
      END
   END n_16680

   PIN n_16684
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.85 187.49 307.95 188 ;
      END
   END n_16684

   PIN n_212558
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 255.85 187.49 255.95 188 ;
      END
   END n_212558

   PIN n_82772
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 131.55 333.2 131.65 ;
      END
   END n_82772

   PIN n_82780
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 135.55 333.2 135.65 ;
      END
   END n_82780

   PIN n_82909
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 146.75 333.2 146.85 ;
      END
   END n_82909

   PIN n_83007
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 130.15 333.2 130.25 ;
      END
   END n_83007

   PIN n_83063
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 35.95 333.2 36.05 ;
      END
   END n_83063

   PIN n_83143
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 127.15 333.2 127.25 ;
      END
   END n_83143

   PIN n_83196
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 147.15 333.2 147.25 ;
      END
   END n_83196

   PIN n_83220
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 151.55 333.2 151.65 ;
      END
   END n_83220

   PIN n_83253
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.945 153.9 333.2 154.1 ;
      END
   END n_83253

   PIN n_83284
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 148.75 333.2 148.85 ;
      END
   END n_83284

   PIN n_83297
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 94.75 333.2 94.85 ;
      END
   END n_83297

   PIN n_83370
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 122.35 333.2 122.45 ;
      END
   END n_83370

   PIN n_83394
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 144.15 333.2 144.25 ;
      END
   END n_83394

   PIN n_83464
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 121.35 333.2 121.45 ;
      END
   END n_83464

   PIN n_83518
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 121.75 333.2 121.85 ;
      END
   END n_83518

   PIN n_83537
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 151.35 333.2 151.45 ;
      END
   END n_83537

   PIN n_83544
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 142.35 333.2 142.45 ;
      END
   END n_83544

   PIN n_83637
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 134.75 333.2 134.85 ;
      END
   END n_83637

   PIN n_83660
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 152.95 333.2 153.05 ;
      END
   END n_83660

   PIN n_83662
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 118.95 333.2 119.05 ;
      END
   END n_83662

   PIN n_83713
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 130.55 333.2 130.65 ;
      END
   END n_83713

   PIN n_83717
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 143.95 333.2 144.05 ;
      END
   END n_83717

   PIN n_83770
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 122.55 333.2 122.65 ;
      END
   END n_83770

   PIN n_83804
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 12.15 333.2 12.25 ;
      END
   END n_83804

   PIN n_83818
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 141.75 333.2 141.85 ;
      END
   END n_83818

   PIN n_83848
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 141.75 333.2 141.85 ;
      END
   END n_83848

   PIN n_83939
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.945 24.3 333.2 24.5 ;
      END
   END n_83939

   PIN n_83944
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 123.15 333.2 123.25 ;
      END
   END n_83944

   PIN n_84141
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 146.55 333.2 146.65 ;
      END
   END n_84141

   PIN n_84142
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 305.05 0 305.15 0.51 ;
      END
   END n_84142

   PIN n_84180
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 127.35 333.2 127.45 ;
      END
   END n_84180

   PIN n_84307
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 280.85 187.49 280.95 188 ;
      END
   END n_84307

   PIN n_84316
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 121.15 333.2 121.25 ;
      END
   END n_84316

   PIN n_84391
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 123.35 333.2 123.45 ;
      END
   END n_84391

   PIN n_84580
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 126.95 333.2 127.05 ;
      END
   END n_84580

   PIN n_84632
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 148.55 333.2 148.65 ;
      END
   END n_84632

   PIN n_84645
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 125.35 333.2 125.45 ;
      END
   END n_84645

   PIN n_84646
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 125.15 333.2 125.25 ;
      END
   END n_84646

   PIN n_84687
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 128.55 333.2 128.65 ;
      END
   END n_84687

   PIN n_84688
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 128.35 333.2 128.45 ;
      END
   END n_84688

   PIN n_84801
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 137.15 333.2 137.25 ;
      END
   END n_84801

   PIN n_84811
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 146.95 333.2 147.05 ;
      END
   END n_84811

   PIN n_84823
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 126.95 333.2 127.05 ;
      END
   END n_84823

   PIN n_84840
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 156.55 333.2 156.65 ;
      END
   END n_84840

   PIN n_84875
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 122.95 333.2 123.05 ;
      END
   END n_84875

   PIN n_84895
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.65 187.49 321.75 188 ;
      END
   END n_84895

   PIN n_84903
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 136.15 333.2 136.25 ;
      END
   END n_84903

   PIN n_84918
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 317.85 187.49 317.95 188 ;
      END
   END n_84918

   PIN n_84940
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 146.35 333.2 146.45 ;
      END
   END n_84940

   PIN n_84990
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.25 187.49 320.35 188 ;
      END
   END n_84990

   PIN n_85014
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 142.95 333.2 143.05 ;
      END
   END n_85014

   PIN n_85057
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 89.05 187.49 89.15 188 ;
      END
   END n_85057

   PIN n_85084
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 142.55 333.2 142.65 ;
      END
   END n_85084

   PIN n_85194
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 168.35 333.2 168.45 ;
      END
   END n_85194

   PIN n_85234
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 268.45 187.49 268.55 188 ;
      END
   END n_85234

   PIN n_85248
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 283.65 187.49 283.75 188 ;
      END
   END n_85248

   PIN n_85335
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.45 187.49 306.55 188 ;
      END
   END n_85335

   PIN n_85437
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.945 147.7 333.2 147.9 ;
      END
   END n_85437

   PIN n_85457
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 280.65 187.49 280.75 188 ;
      END
   END n_85457

   PIN n_85462
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.45 187.49 293.55 188 ;
      END
   END n_85462

   PIN n_85470
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.65 187.49 320.75 188 ;
      END
   END n_85470

   PIN n_85495
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 317.05 187.49 317.15 188 ;
      END
   END n_85495

   PIN n_85591
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.25 187.49 232.35 188 ;
      END
   END n_85591

   PIN n_85698
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 114.95 333.2 115.05 ;
      END
   END n_85698

   PIN n_85825
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 280.45 187.49 280.55 188 ;
      END
   END n_85825

   PIN n_85840
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 268.25 187.49 268.35 188 ;
      END
   END n_85840

   PIN n_85969
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 280.25 187.49 280.35 188 ;
      END
   END n_85969

   PIN n_85975
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 268.05 187.49 268.15 188 ;
      END
   END n_85975

   PIN n_86111
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.85 187.49 267.95 188 ;
      END
   END n_86111

   PIN n_86144
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 156.15 333.2 156.25 ;
      END
   END n_86144

   PIN n_86164
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 171.15 333.2 171.25 ;
      END
   END n_86164

   PIN n_86241
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 280.05 187.49 280.15 188 ;
      END
   END n_86241

   PIN n_86242
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.85 187.49 244.95 188 ;
      END
   END n_86242

   PIN n_86243
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.25 187.49 293.35 188 ;
      END
   END n_86243

   PIN n_86295
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 169.55 333.2 169.65 ;
      END
   END n_86295

   PIN n_86457
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 169.35 333.2 169.45 ;
      END
   END n_86457

   PIN n_86466
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 155.75 333.2 155.85 ;
      END
   END n_86466

   PIN n_86468
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 179.95 333.2 180.05 ;
      END
   END n_86468

   PIN n_86472
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 290.65 187.49 290.75 188 ;
      END
   END n_86472

   PIN n_86473
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 290.45 187.49 290.55 188 ;
      END
   END n_86473

   PIN n_86493
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.65 187.49 270.75 188 ;
      END
   END n_86493

   PIN n_86500
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.65 187.49 267.75 188 ;
      END
   END n_86500

   PIN n_86542
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 169.15 333.2 169.25 ;
      END
   END n_86542

   PIN n_86577
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 170.95 333.2 171.05 ;
      END
   END n_86577

   PIN n_86583
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 295.25 187.49 295.35 188 ;
      END
   END n_86583

   PIN n_86594
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 305.65 187.49 305.75 188 ;
      END
   END n_86594

   PIN n_86596
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.85 187.49 279.95 188 ;
      END
   END n_86596

   PIN n_86598
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 280.45 187.49 280.55 188 ;
      END
   END n_86598

   PIN n_86602
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 152.75 333.2 152.85 ;
      END
   END n_86602

   PIN n_86605
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.45 187.49 267.55 188 ;
      END
   END n_86605

   PIN n_86618
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 170.75 333.2 170.85 ;
      END
   END n_86618

   PIN n_86641
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 267.65 187.49 267.75 188 ;
      END
   END n_86641

   PIN n_86642
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 154.55 333.2 154.65 ;
      END
   END n_86642

   PIN n_86644
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 267.45 187.49 267.55 188 ;
      END
   END n_86644

   PIN n_86648
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 141.15 333.2 141.25 ;
      END
   END n_86648

   PIN n_86690
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 304.25 187.49 304.35 188 ;
      END
   END n_86690

   PIN n_86691
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.65 187.49 291.75 188 ;
      END
   END n_86691

   PIN n_86696
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 133.95 333.2 134.05 ;
      END
   END n_86696

   PIN n_86750
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 290.25 187.49 290.35 188 ;
      END
   END n_86750

   PIN n_86804
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.65 187.49 279.75 188 ;
      END
   END n_86804

   PIN n_86806
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.25 187.49 267.35 188 ;
      END
   END n_86806

   PIN n_86807
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.45 187.49 291.55 188 ;
      END
   END n_86807

   PIN n_86815
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.85 187.49 320.95 188 ;
      END
   END n_86815

   PIN n_86816
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 321.05 187.49 321.15 188 ;
      END
   END n_86816

   PIN n_86829
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 279.45 187.49 279.55 188 ;
      END
   END n_86829

   PIN n_86839
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 301.45 187.49 301.55 188 ;
      END
   END n_86839

   PIN n_86843
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 143.75 333.2 143.85 ;
      END
   END n_86843

   PIN n_86851
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 181.55 333.2 181.65 ;
      END
   END n_86851

   PIN n_86861
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 116.35 333.2 116.45 ;
      END
   END n_86861

   PIN n_86969
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.45 187.49 234.55 188 ;
      END
   END n_86969

   PIN n_87008
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 134.95 333.2 135.05 ;
      END
   END n_87008

   PIN n_87034
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.05 187.49 234.15 188 ;
      END
   END n_87034

   PIN n_87060
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 85.95 333.2 86.05 ;
      END
   END n_87060

   PIN n_87145
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 102.95 333.2 103.05 ;
      END
   END n_87145

   PIN n_87155
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 90.95 333.2 91.05 ;
      END
   END n_87155

   PIN n_87159
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 96.95 333.2 97.05 ;
      END
   END n_87159

   PIN n_87178
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 293.25 187.49 293.35 188 ;
      END
   END n_87178

   PIN n_87180
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 245.65 187.49 245.75 188 ;
      END
   END n_87180

   PIN n_87185
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 154.55 333.2 154.65 ;
      END
   END n_87185

   PIN n_87213
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 131.35 333.2 131.45 ;
      END
   END n_87213

   PIN n_87230
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 285.45 187.49 285.55 188 ;
      END
   END n_87230

   PIN n_87235
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 157.55 333.2 157.65 ;
      END
   END n_87235

   PIN n_87275
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 147.55 333.2 147.65 ;
      END
   END n_87275

   PIN n_87293
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 258.05 187.49 258.15 188 ;
      END
   END n_87293

   PIN n_87322
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.65 187.49 244.75 188 ;
      END
   END n_87322

   PIN n_87328
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 97.95 333.2 98.05 ;
      END
   END n_87328

   PIN n_87329
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 95.55 333.2 95.65 ;
      END
   END n_87329

   PIN n_87354
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 305.25 187.49 305.35 188 ;
      END
   END n_87354

   PIN n_87367
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 221.85 187.49 221.95 188 ;
      END
   END n_87367

   PIN n_87409
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.45 187.49 244.55 188 ;
      END
   END n_87409

   PIN n_87410
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.25 187.49 244.35 188 ;
      END
   END n_87410

   PIN n_87427
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.05 187.49 306.15 188 ;
      END
   END n_87427

   PIN n_87453
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.45 187.49 294.55 188 ;
      END
   END n_87453

   PIN n_87468
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 246.45 187.49 246.55 188 ;
      END
   END n_87468

   PIN n_87487
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 234 187.745 234.2 188 ;
      END
   END n_87487

   PIN n_87488
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 267.05 187.49 267.15 188 ;
      END
   END n_87488

   PIN n_87493
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 92.95 333.2 93.05 ;
      END
   END n_87493

   PIN n_87500
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 247.05 187.49 247.15 188 ;
      END
   END n_87500

   PIN n_87508
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.45 187.49 245.55 188 ;
      END
   END n_87508

   PIN n_87509
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 244.05 187.49 244.15 188 ;
      END
   END n_87509

   PIN n_87518
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 268.85 187.49 268.95 188 ;
      END
   END n_87518

   PIN n_87532
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 246.25 187.49 246.35 188 ;
      END
   END n_87532

   PIN n_87574
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.65 187.49 220.75 188 ;
      END
   END n_87574

   PIN n_87595
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 151.15 333.2 151.25 ;
      END
   END n_87595

   PIN n_87624
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.85 187.49 266.95 188 ;
      END
   END n_87624

   PIN n_87630
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 232.05 187.49 232.15 188 ;
      END
   END n_87630

   PIN n_87656
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 246.05 187.49 246.15 188 ;
      END
   END n_87656

   PIN n_87658
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 294.25 187.49 294.35 188 ;
      END
   END n_87658

   PIN n_87663
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.85 187.49 257.95 188 ;
      END
   END n_87663

   PIN n_87665
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 305.05 187.49 305.15 188 ;
      END
   END n_87665

   PIN n_87666
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 255.05 187.49 255.15 188 ;
      END
   END n_87666

   PIN n_87668
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 98.95 333.2 99.05 ;
      END
   END n_87668

   PIN n_87689
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 148.35 333.2 148.45 ;
      END
   END n_87689

   PIN n_87742
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.85 187.49 233.95 188 ;
      END
   END n_87742

   PIN n_87751
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 245.45 187.49 245.55 188 ;
      END
   END n_87751

   PIN n_87756
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 305.85 187.49 305.95 188 ;
      END
   END n_87756

   PIN n_87776
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 152.55 333.2 152.65 ;
      END
   END n_87776

   PIN n_87779
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.25 187.49 245.35 188 ;
      END
   END n_87779

   PIN n_87782
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 243.85 187.49 243.95 188 ;
      END
   END n_87782

   PIN n_87803
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 97.55 333.2 97.65 ;
      END
   END n_87803

   PIN n_87807
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 208.85 187.49 208.95 188 ;
      END
   END n_87807

   PIN n_87810
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.45 187.49 220.55 188 ;
      END
   END n_87810

   PIN n_87819
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 231.85 187.49 231.95 188 ;
      END
   END n_87819

   PIN n_87842
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 152.35 333.2 152.45 ;
      END
   END n_87842

   PIN n_87860
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.25 187.49 220.35 188 ;
      END
   END n_87860

   PIN n_87863
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 257.25 187.49 257.35 188 ;
      END
   END n_87863

   PIN n_87872
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.65 187.49 266.75 188 ;
      END
   END n_87872

   PIN n_87884
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 231.85 187.49 231.95 188 ;
      END
   END n_87884

   PIN n_87897
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 196.45 187.49 196.55 188 ;
      END
   END n_87897

   PIN n_87911
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 136.35 333.2 136.45 ;
      END
   END n_87911

   PIN n_87937
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 125.05 187.49 125.15 188 ;
      END
   END n_87937

   PIN n_87953
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 157.35 333.2 157.45 ;
      END
   END n_87953

   PIN n_87954
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 143.55 333.2 143.65 ;
      END
   END n_87954

   PIN n_87964
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.25 187.49 306.35 188 ;
      END
   END n_87964

   PIN n_87971
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 68.95 333.2 69.05 ;
      END
   END n_87971

   PIN n_87976
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 100.95 333.2 101.05 ;
      END
   END n_87976

   PIN n_87986
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.45 187.49 279.55 188 ;
      END
   END n_87986

   PIN n_88058
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 293.05 187.49 293.15 188 ;
      END
   END n_88058

   PIN n_88113
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 231.65 187.49 231.75 188 ;
      END
   END n_88113

   PIN n_88117
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 83.75 333.2 83.85 ;
      END
   END n_88117

   PIN n_88193
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 138.35 333.2 138.45 ;
      END
   END n_88193

   PIN n_88207
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 245.25 187.49 245.35 188 ;
      END
   END n_88207

   PIN n_88213
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 154.75 333.2 154.85 ;
      END
   END n_88213

   PIN n_88245
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 266.45 187.49 266.55 188 ;
      END
   END n_88245

   PIN n_88254
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 141.55 333.2 141.65 ;
      END
   END n_88254

   PIN n_88256
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.85 187.49 318.95 188 ;
      END
   END n_88256

   PIN n_88259
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.05 187.49 319.15 188 ;
      END
   END n_88259

   PIN n_88261
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.25 187.49 291.35 188 ;
      END
   END n_88261

   PIN n_88265
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 137.95 333.2 138.05 ;
      END
   END n_88265

   PIN n_88318
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 150.95 333.2 151.05 ;
      END
   END n_88318

   PIN n_88320
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 129.75 333.2 129.85 ;
      END
   END n_88320

   PIN n_88346
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 143.35 333.2 143.45 ;
      END
   END n_88346

   PIN n_88381
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 220.05 187.49 220.15 188 ;
      END
   END n_88381

   PIN n_88397
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 143.15 333.2 143.25 ;
      END
   END n_88397

   PIN n_88416
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 291.05 187.49 291.15 188 ;
      END
   END n_88416

   PIN n_88417
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 290.85 187.49 290.95 188 ;
      END
   END n_88417

   PIN n_88426
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 152.15 333.2 152.25 ;
      END
   END n_88426

   PIN n_88428
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 155.95 333.2 156.05 ;
      END
   END n_88428

   PIN n_88454
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 153.55 333.2 153.65 ;
      END
   END n_88454

   PIN n_88468
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 172.85 187.49 172.95 188 ;
      END
   END n_88468

   PIN n_88469
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 290.65 187.49 290.75 188 ;
      END
   END n_88469

   PIN n_88523
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 234.25 187.49 234.35 188 ;
      END
   END n_88523

   PIN n_88555
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 141.35 333.2 141.45 ;
      END
   END n_88555

   PIN n_88572
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 231.65 187.49 231.75 188 ;
      END
   END n_88572

   PIN n_88589
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 290.45 187.49 290.55 188 ;
      END
   END n_88589

   PIN n_88594
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 243.65 187.49 243.75 188 ;
      END
   END n_88594

   PIN n_88626
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 157.15 333.2 157.25 ;
      END
   END n_88626

   PIN n_88646
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 131.75 333.2 131.85 ;
      END
   END n_88646

   PIN n_88652
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 246.85 187.49 246.95 188 ;
      END
   END n_88652

   PIN n_88668
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 155.75 333.2 155.85 ;
      END
   END n_88668

   PIN n_88683
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 290.25 187.49 290.35 188 ;
      END
   END n_88683

   PIN n_88697
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 255.65 187.49 255.75 188 ;
      END
   END n_88697

   PIN n_88703
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 306.65 187.49 306.75 188 ;
      END
   END n_88703

   PIN n_88704
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 255.45 187.49 255.55 188 ;
      END
   END n_88704

   PIN n_88705
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.25 187.49 279.35 188 ;
      END
   END n_88705

   PIN n_88706
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 243.45 187.49 243.55 188 ;
      END
   END n_88706

   PIN n_88707
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 279.05 187.49 279.15 188 ;
      END
   END n_88707

   PIN n_88708
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 278.85 187.49 278.95 188 ;
      END
   END n_88708

   PIN n_88786
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.45 187.49 270.55 188 ;
      END
   END n_88786

   PIN n_88805
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 279.25 187.49 279.35 188 ;
      END
   END n_88805

   PIN n_88833
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 124.95 333.2 125.05 ;
      END
   END n_88833

   PIN n_88835
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 267.25 187.49 267.35 188 ;
      END
   END n_88835

   PIN n_88854
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 127.15 333.2 127.25 ;
      END
   END n_88854

   PIN n_89083
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 267.05 187.49 267.15 188 ;
      END
   END n_89083

   PIN n_89164
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 266.85 187.49 266.95 188 ;
      END
   END n_89164

   PIN n_89232
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 312.45 187.49 312.55 188 ;
      END
   END n_89232

   PIN n_89272
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 313.85 187.49 313.95 188 ;
      END
   END n_89272

   PIN n_89334
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 316.65 187.49 316.75 188 ;
      END
   END n_89334

   PIN n_89338
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 312.65 187.49 312.75 188 ;
      END
   END n_89338

   PIN n_89339
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 317.25 187.49 317.35 188 ;
      END
   END n_89339

   PIN n_89351
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 310.05 187.49 310.15 188 ;
      END
   END n_89351

   PIN n_89410
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 308.6 187.745 308.8 188 ;
      END
   END n_89410

   PIN n_89426
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 311.45 187.49 311.55 188 ;
      END
   END n_89426

   PIN n_89435
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 310.45 187.49 310.55 188 ;
      END
   END n_89435

   PIN n_89436
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 294.25 187.49 294.35 188 ;
      END
   END n_89436

   PIN n_89496
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 312.85 187.49 312.95 188 ;
      END
   END n_89496

   PIN n_89517
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 311.65 187.49 311.75 188 ;
      END
   END n_89517

   PIN n_89518
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 309.65 187.49 309.75 188 ;
      END
   END n_89518

   PIN n_89528
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 318.45 187.49 318.55 188 ;
      END
   END n_89528

   PIN n_89581
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 310.25 187.49 310.35 188 ;
      END
   END n_89581

   PIN n_89657
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 309.65 187.49 309.75 188 ;
      END
   END n_89657

   PIN n_89673
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 314.65 187.49 314.75 188 ;
      END
   END n_89673

   PIN n_89840
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 307.05 187.49 307.15 188 ;
      END
   END n_89840

   PIN n_89892
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 149.75 333.2 149.85 ;
      END
   END n_89892

   PIN n_89963
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 311.45 187.49 311.55 188 ;
      END
   END n_89963

   PIN n_90020
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 140.35 333.2 140.45 ;
      END
   END n_90020

   PIN n_90052
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 311.25 187.49 311.35 188 ;
      END
   END n_90052

   PIN n_90172
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 292.85 187.49 292.95 188 ;
      END
   END n_90172

   PIN n_90334
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 231.45 187.49 231.55 188 ;
      END
   END n_90334

   PIN n_90504
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 307.25 187.49 307.35 188 ;
      END
   END n_90504

   PIN n_90645
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 312.85 187.49 312.95 188 ;
      END
   END n_90645

   PIN n_90656
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 208.65 187.49 208.75 188 ;
      END
   END n_90656

   PIN n_90669
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 148.15 333.2 148.25 ;
      END
   END n_90669

   PIN n_90684
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 147.95 333.2 148.05 ;
      END
   END n_90684

   PIN n_90710
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.25 187.49 270.35 188 ;
      END
   END n_90710

   PIN n_90712
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 146.15 333.2 146.25 ;
      END
   END n_90712

   PIN u2_L2_reg_17__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 129.55 333.2 129.65 ;
      END
   END u2_L2_reg_17__Q

   PIN u2_L2_reg_9__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 127.35 333.2 127.45 ;
      END
   END u2_L2_reg_9__Q

   PIN u2_L3_reg_17__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 140.95 333.2 141.05 ;
      END
   END u2_L3_reg_17__Q

   PIN u2_L3_reg_9__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 309.25 187.49 309.35 188 ;
      END
   END u2_L3_reg_9__Q

   PIN u2_L4_12_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 110.95 333.2 111.05 ;
      END
   END u2_L4_12_

   PIN u2_L4_19_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 231.25 187.49 231.35 188 ;
      END
   END u2_L4_19_

   PIN u2_L4_22_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 318.65 187.49 318.75 188 ;
      END
   END u2_L4_22_

   PIN u2_L4_29_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 106.95 333.2 107.05 ;
      END
   END u2_L4_29_

   PIN u2_L4_reg_7__Q
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 103.15 333.2 103.25 ;
      END
   END u2_L4_reg_7__Q

   PIN u2_R2_13_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 123.75 333.2 123.85 ;
      END
   END u2_R2_13_

   PIN u2_R2_14_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 136.95 333.2 137.05 ;
      END
   END u2_R2_14_

   PIN u2_R2_28_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 116.95 333.2 117.05 ;
      END
   END u2_R2_28_

   PIN u2_R2_2_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 142.95 333.2 143.05 ;
      END
   END u2_R2_2_

   PIN u2_R3_11_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 134.35 333.2 134.45 ;
      END
   END u2_R3_11_

   PIN u2_R3_12_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 129.35 333.2 129.45 ;
      END
   END u2_R3_12_

   PIN u2_R3_17_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 129.15 333.2 129.25 ;
      END
   END u2_R3_17_

   PIN u2_R3_18_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 135.55 333.2 135.65 ;
      END
   END u2_R3_18_

   PIN u2_R3_22_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 155.55 333.2 155.65 ;
      END
   END u2_R3_22_

   PIN u2_R3_23_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 131.35 333.2 131.45 ;
      END
   END u2_R3_23_

   PIN u2_R3_26_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 305.05 0 305.15 0.51 ;
      END
   END u2_R3_26_

   PIN u2_R3_28_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 135.75 333.2 135.85 ;
      END
   END u2_R3_28_

   PIN u2_R3_31_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 140.95 333.2 141.05 ;
      END
   END u2_R3_31_

   PIN u2_R3_3_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 307.65 187.49 307.75 188 ;
      END
   END u2_R3_3_

   PIN u2_R3_4_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 131.15 333.2 131.25 ;
      END
   END u2_R3_4_

   PIN u2_R3_5_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 322.25 187.49 322.35 188 ;
      END
   END u2_R3_5_

   PIN u2_R3_8_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 130.35 333.2 130.45 ;
      END
   END u2_R3_8_

   PIN u2_R4_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 332.69 149.55 333.2 149.65 ;
      END
   END u2_R4_10_

   PIN u2_R4_12_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 140.15 333.2 140.25 ;
      END
   END u2_R4_12_

   PIN u2_R4_14_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 320.05 187.49 320.15 188 ;
      END
   END u2_R4_14_

   PIN u2_R4_24_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 245.85 187.49 245.95 188 ;
      END
   END u2_R4_24_

   PIN u2_R4_26_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 320.45 187.49 320.55 188 ;
      END
   END u2_R4_26_

   PIN u2_R4_30_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 317.25 187.49 317.35 188 ;
      END
   END u2_R4_30_

   PIN u2_R4_31_
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 332.69 131.15 333.2 131.25 ;
      END
   END u2_R4_31_

   PIN u2_uk_K_r_420
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 319.25 187.49 319.35 188 ;
      END
   END u2_uk_K_r_420

   OBS
      LAYER via4 ;
         RECT 0 0 333.2 188 ;
      LAYER via1 ;
         RECT 0 0 333.2 188 ;
      LAYER metal5 ;
         RECT 0 0 333.2 188 ;
      LAYER metal4 ;
         RECT 0 0 333.2 188 ;
      LAYER metal3 ;
         RECT 0 0 333.2 188 ;
      LAYER metal2 ;
         RECT 0 0 333.2 188 ;
      LAYER metal1 ;
         RECT 0 0 333.2 188 ;
   END
END h1

MACRO h0
   CLASS BLOCK ;
   FOREIGN h0 ;
   ORIGIN 0 0 ;
   SIZE 280 BY 296.81 ;
   SYMMETRY X Y R90 ;
   PIN FE_OFN2124_n_92148
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 135.35 280 135.45 ;
      END
   END FE_OFN2124_n_92148

   PIN FE_OFN2215_n_2854
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 119.85 0 119.95 0.51 ;
      END
   END FE_OFN2215_n_2854

   PIN g202734_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 148.15 280 148.25 ;
      END
   END g202734_p

   PIN g289278_p2
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.85 0 91.95 0.51 ;
      END
   END g289278_p2

   PIN g289637_p1
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.05 0 151.15 0.51 ;
      END
   END g289637_p1

   PIN g291339_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 132.05 0 132.15 0.51 ;
      END
   END g291339_p

   PIN g301491_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.75 0.51 39.85 ;
      END
   END g301491_p

   PIN g302166_p
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 71.15 0.51 71.25 ;
      END
   END g302166_p

   PIN key_c_r_26__2568
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 87.25 0 87.35 0.51 ;
      END
   END key_c_r_26__2568

   PIN n_10300
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.65 0 115.75 0.51 ;
      END
   END n_10300

   PIN n_10543
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.25 0 138.35 0.51 ;
      END
   END n_10543

   PIN n_10664
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.05 0 141.15 0.51 ;
      END
   END n_10664

   PIN n_11092
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 139.85 0 139.95 0.51 ;
      END
   END n_11092

   PIN n_11160
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.65 0 116.75 0.51 ;
      END
   END n_11160

   PIN n_11190
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 129.85 0 129.95 0.51 ;
      END
   END n_11190

   PIN n_11283
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.85 0 115.95 0.51 ;
      END
   END n_11283

   PIN n_116769
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.65 0 199.75 0.51 ;
      END
   END n_116769

   PIN n_116784
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.25 0 20.35 0.51 ;
      END
   END n_116784

   PIN n_117640
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.85 0 141.95 0.51 ;
      END
   END n_117640

   PIN n_117987
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 191.85 0 191.95 0.51 ;
      END
   END n_117987

   PIN n_1204
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 202.65 0 202.75 0.51 ;
      END
   END n_1204

   PIN n_1209
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 172.15 0.51 172.25 ;
      END
   END n_1209

   PIN n_12805
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.05 0 80.15 0.51 ;
      END
   END n_12805

   PIN n_12937
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 96.05 0 96.15 0.51 ;
      END
   END n_12937

   PIN n_12977
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 79.85 0 79.95 0.51 ;
      END
   END n_12977

   PIN n_1417
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 186.85 0 186.95 0.51 ;
      END
   END n_1417

   PIN n_14736
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 226.05 0 226.15 0.51 ;
      END
   END n_14736

   PIN n_1579
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 205.85 0 205.95 0.51 ;
      END
   END n_1579

   PIN n_17638
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 228.45 0 228.55 0.51 ;
      END
   END n_17638

   PIN n_18022
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.05 0 272.15 0.51 ;
      END
   END n_18022

   PIN n_18160
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 15.55 280 15.65 ;
      END
   END n_18160

   PIN n_2208
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.35 0.51 28.45 ;
      END
   END n_2208

   PIN n_2598
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.15 0.51 52.25 ;
      END
   END n_2598

   PIN n_3390
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 52.15 0.51 52.25 ;
      END
   END n_3390

   PIN n_3453
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 39.95 0.51 40.05 ;
      END
   END n_3453

   PIN n_3518
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.05 0 92.15 0.51 ;
      END
   END n_3518

   PIN n_3653
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.35 0.51 40.45 ;
      END
   END n_3653

   PIN n_3919
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 82.95 0.51 83.05 ;
      END
   END n_3919

   PIN n_4023
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.85 0 67.95 0.51 ;
      END
   END n_4023

   PIN n_4025
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 63.95 0.51 64.05 ;
      END
   END n_4025

   PIN n_4166
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 68.05 0 68.15 0.51 ;
      END
   END n_4166

   PIN n_4717
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 64.15 0.51 64.25 ;
      END
   END n_4717

   PIN n_4718
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.75 0.51 52.85 ;
      END
   END n_4718

   PIN n_4927
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.35 0.51 52.45 ;
      END
   END n_4927

   PIN n_5717
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 112.15 0.51 112.25 ;
      END
   END n_5717

   PIN n_66187
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 64.15 280 64.25 ;
      END
   END n_66187

   PIN n_66261
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 64.35 280 64.45 ;
      END
   END n_66261

   PIN n_7078
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 236.25 0 236.35 0.51 ;
      END
   END n_7078

   PIN n_7087
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 143.85 0 143.95 0.51 ;
      END
   END n_7087

   PIN n_7431
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 211.45 0 211.55 0.51 ;
      END
   END n_7431

   PIN n_7877
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 158.85 0 158.95 0.51 ;
      END
   END n_7877

   PIN n_8063
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.65 0 140.75 0.51 ;
      END
   END n_8063

   PIN n_8726
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 156.25 0 156.35 0.51 ;
      END
   END n_8726

   PIN n_8829
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 157.65 0 157.75 0.51 ;
      END
   END n_8829

   PIN n_91001
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 123.95 280 124.05 ;
      END
   END n_91001

   PIN n_9103
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 154.85 0 154.95 0.51 ;
      END
   END n_9103

   PIN n_91121
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 87.95 280 88.05 ;
      END
   END n_91121

   PIN n_91266
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 28.15 280 28.25 ;
      END
   END n_91266

   PIN n_91489
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 28.75 280 28.85 ;
      END
   END n_91489

   PIN n_91525
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 100.35 280 100.45 ;
      END
   END n_91525

   PIN n_91573
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 15.75 280 15.85 ;
      END
   END n_91573

   PIN n_91692
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 99.75 280 99.85 ;
      END
   END n_91692

   PIN n_91814
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 100.55 280 100.65 ;
      END
   END n_91814

   PIN n_91815
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 13.75 280 13.85 ;
      END
   END n_91815

   PIN n_91824
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 124.35 280 124.45 ;
      END
   END n_91824

   PIN n_91825
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 135.95 280 136.05 ;
      END
   END n_91825

   PIN n_91826
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 99.95 280 100.05 ;
      END
   END n_91826

   PIN n_91828
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 112.15 280 112.25 ;
      END
   END n_91828

   PIN n_91839
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 112.35 280 112.45 ;
      END
   END n_91839

   PIN n_91845
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 28.35 280 28.45 ;
      END
   END n_91845

   PIN n_92019
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 27.95 280 28.05 ;
      END
   END n_92019

   PIN n_92117
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 112.55 280 112.65 ;
      END
   END n_92117

   PIN n_92305
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 15.95 280 16.05 ;
      END
   END n_92305

   PIN n_92419
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 112.75 280 112.85 ;
      END
   END n_92419

   PIN n_92502
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal5 ;
             RECT 279.49 11.75 280 11.85 ;
      END
   END n_92502

   PIN n_92510
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 28.55 280 28.65 ;
      END
   END n_92510

   PIN n_92511
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 136.15 280 136.25 ;
      END
   END n_92511

   PIN n_9282
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.65 0 159.75 0.51 ;
      END
   END n_9282

   PIN n_95488
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 148.35 280 148.45 ;
      END
   END n_95488

   PIN n_95562
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 16.15 280 16.25 ;
      END
   END n_95562

   PIN n_95579
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 12.15 280 12.25 ;
      END
   END n_95579

   PIN n_95580
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 148.55 280 148.65 ;
      END
   END n_95580

   PIN n_95719
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 160.15 280 160.25 ;
      END
   END n_95719

   PIN n_95756
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 28.95 280 29.05 ;
      END
   END n_95756

   PIN n_95826
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.745 11.1 280 11.3 ;
      END
   END n_95826

   PIN n_95913
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 172.15 280 172.25 ;
      END
   END n_95913

   PIN n_95976
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 29.15 280 29.25 ;
      END
   END n_95976

   PIN n_96109
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 148.75 280 148.85 ;
      END
   END n_96109

   PIN n_96227
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 160.35 280 160.45 ;
      END
   END n_96227

   PIN n_96448
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 29.35 280 29.45 ;
      END
   END n_96448

   PIN n_96488
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 40.15 280 40.25 ;
      END
   END n_96488

   PIN n_9734
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 156.65 0 156.75 0.51 ;
      END
   END n_9734

   PIN u0_L0_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.45 0 8.55 0.51 ;
      END
   END u0_L0_10_

   PIN u0_L0_4_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.25 0 80.35 0.51 ;
      END
   END u0_L0_4_

   PIN u0_L0_6_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 140.05 0 140.15 0.51 ;
      END
   END u0_L0_6_

   PIN u0_L1_10_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 229.45 0 229.55 0.51 ;
      END
   END u0_L1_10_

   PIN u0_L1_1_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 175.85 0 175.95 0.51 ;
      END
   END u0_L1_1_

   PIN u0_R0_23_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 109.05 0 109.15 0.51 ;
      END
   END u0_R0_23_

   PIN u0_R0_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal4 ;
             RECT 184.65 0 184.75 0.51 ;
      END
   END u0_R0_28_

   PIN u1_key_r_28_
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 133.35 280 133.45 ;
      END
   END u1_key_r_28_

   PIN FE_OFN1268_n_3950
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 88.95 0.51 89.05 ;
      END
   END FE_OFN1268_n_3950

   PIN FE_OFN1270_n_6370
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 100.15 0.51 100.25 ;
      END
   END FE_OFN1270_n_6370

   PIN FE_OFN1342_n_5733
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 111.05 0 111.15 0.51 ;
      END
   END FE_OFN1342_n_5733

   PIN FE_OFN1346_n_1012
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 188.05 0 188.15 0.51 ;
      END
   END FE_OFN1346_n_1012

   PIN FE_OFN1882_n_1371
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 83.95 0.51 84.05 ;
      END
   END FE_OFN1882_n_1371

   PIN FE_OFN2123_n_92148
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 88.35 280 88.45 ;
      END
   END FE_OFN2123_n_92148

   PIN FE_OFN2356_n_1288
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 145.45 0 145.55 0.51 ;
      END
   END FE_OFN2356_n_1288

   PIN FE_OFN749_n_15670
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 199.85 0 199.95 0.51 ;
      END
   END FE_OFN749_n_15670

   PIN desIn_13_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 16.15 0.51 16.25 ;
      END
   END desIn_13_

   PIN desIn_31_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 15.95 0.51 16.05 ;
      END
   END desIn_31_

   PIN desIn_38_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.05 296.2961 272.15 296.8061 ;
      END
   END desIn_38_

   PIN desIn_50_
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 40.15 0.51 40.25 ;
      END
   END desIn_50_

   PIN g303844_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 248.05 0 248.15 0.51 ;
      END
   END g303844_db

   PIN g303844_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.05 0 260.15 0.51 ;
      END
   END g303844_sb

   PIN g321474_db
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.25 0 8.35 0.51 ;
      END
   END g321474_db

   PIN g321474_sb
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 70.85 0 70.95 0.51 ;
      END
   END g321474_sb

   PIN ispd_clk
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.745 132.9 280 133.1 ;
      END
   END ispd_clk

   PIN key_b_r_16__28_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 80.05 296.2961 80.15 296.8061 ;
      END
   END key_b_r_16__28_

   PIN key_c_r_25__2513
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 88.25 296.2961 88.35 296.8061 ;
      END
   END key_c_r_25__2513

   PIN n_10016
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.85 0 103.95 0.51 ;
      END
   END n_10016

   PIN n_10047
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.45 0 116.55 0.51 ;
      END
   END n_10047

   PIN n_10087
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 129.25 0 129.35 0.51 ;
      END
   END n_10087

   PIN n_10299
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 138.65 0 138.75 0.51 ;
      END
   END n_10299

   PIN n_10307
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 104.05 0 104.15 0.51 ;
      END
   END n_10307

   PIN n_10322
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 128.05 0 128.15 0.51 ;
      END
   END n_10322

   PIN n_10332
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 116.2 0 116.4 0.255 ;
      END
   END n_10332

   PIN n_10534
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 133.05 0 133.15 0.51 ;
      END
   END n_10534

   PIN n_10560
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 103.65 0 103.75 0.51 ;
      END
   END n_10560

   PIN n_10579
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 151.45 0 151.55 0.51 ;
      END
   END n_10579

   PIN n_10628
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 129.4 0 129.6 0.255 ;
      END
   END n_10628

   PIN n_10707
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 156.45 0 156.55 0.51 ;
      END
   END n_10707

   PIN n_10905
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 135.45 0 135.55 0.51 ;
      END
   END n_10905

   PIN n_116767
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 218.25 0 218.35 0.51 ;
      END
   END n_116767

   PIN n_116774
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 228.65 0 228.75 0.51 ;
      END
   END n_116774

   PIN n_117986
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 195.45 0 195.55 0.51 ;
      END
   END n_117986

   PIN n_11904
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 131.65 0 131.75 0.51 ;
      END
   END n_11904

   PIN n_11922
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 141.65 0 141.75 0.51 ;
      END
   END n_11922

   PIN n_12137
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.45 0 115.55 0.51 ;
      END
   END n_12137

   PIN n_1241
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 92.25 0 92.35 0.51 ;
      END
   END n_1241

   PIN n_12565
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 91.65 0 91.75 0.51 ;
      END
   END n_12565

   PIN n_1323
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 233.25 0 233.35 0.51 ;
      END
   END n_1323

   PIN n_14285
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 226.25 0 226.35 0.51 ;
      END
   END n_14285

   PIN n_15830
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 176.05 0 176.15 0.51 ;
      END
   END n_15830

   PIN n_15918
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 176.05 0 176.15 0.51 ;
      END
   END n_15918

   PIN n_16285
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 214.65 0 214.75 0.51 ;
      END
   END n_16285

   PIN n_16293
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 188 0 188.2 0.255 ;
      END
   END n_16293

   PIN n_16596
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 220.45 0 220.55 0.51 ;
      END
   END n_16596

   PIN n_16597
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 222.25 0 222.35 0.51 ;
      END
   END n_16597

   PIN n_16611
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 199.85 0 199.95 0.51 ;
      END
   END n_16611

   PIN n_1662
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.15 0.51 77.25 ;
      END
   END n_1662

   PIN n_16731
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 187.65 0 187.75 0.51 ;
      END
   END n_16731

   PIN n_16854
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 218.65 0 218.75 0.51 ;
      END
   END n_16854

   PIN n_1686
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 76.95 0.51 77.05 ;
      END
   END n_1686

   PIN n_16882
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 187.65 0 187.75 0.51 ;
      END
   END n_16882

   PIN n_17069
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 221.85 0 221.95 0.51 ;
      END
   END n_17069

   PIN n_17155
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 216.05 0 216.15 0.51 ;
      END
   END n_17155

   PIN n_1844
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 74.95 0.51 75.05 ;
      END
   END n_1844

   PIN n_1916
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 8.05 0 8.15 0.51 ;
      END
   END n_1916

   PIN n_2108
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 70.95 0.51 71.05 ;
      END
   END n_2108

   PIN n_2210
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.45 0 20.55 0.51 ;
      END
   END n_2210

   PIN n_2597
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 56.05 0 56.15 0.51 ;
      END
   END n_2597

   PIN n_2610
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 8.05 0 8.15 0.51 ;
      END
   END n_2610

   PIN n_2611
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 260.25 0 260.35 0.51 ;
      END
   END n_2611

   PIN n_2721
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 28.15 0.51 28.25 ;
      END
   END n_2721

   PIN n_2854
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 32.05 0 32.15 0.51 ;
      END
   END n_2854

   PIN n_2883
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.95 0.51 52.05 ;
      END
   END n_2883

   PIN n_2885
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 74.3 0.255 74.5 ;
      END
   END n_2885

   PIN n_3058
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 20.05 0 20.15 0.51 ;
      END
   END n_3058

   PIN n_3098
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.75 0.51 51.85 ;
      END
   END n_3098

   PIN n_3175
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.35 0.51 64.45 ;
      END
   END n_3175

   PIN n_3238
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 52.55 0.51 52.65 ;
      END
   END n_3238

   PIN n_3397
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 77.35 0.51 77.45 ;
      END
   END n_3397

   PIN n_3431
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 64.15 0.51 64.25 ;
      END
   END n_3431

   PIN n_3517
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 40.15 0.51 40.25 ;
      END
   END n_3517

   PIN n_3652
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.55 0.51 51.65 ;
      END
   END n_3652

   PIN n_3798
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 89.15 0.51 89.25 ;
      END
   END n_3798

   PIN n_3856
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 27.95 0.51 28.05 ;
      END
   END n_3856

   PIN n_3942
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 80.95 0.51 81.05 ;
      END
   END n_3942

   PIN n_3949
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 99.95 0.51 100.05 ;
      END
   END n_3949

   PIN n_4410
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 51.35 0.51 51.45 ;
      END
   END n_4410

   PIN n_4867
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 100.35 0.51 100.45 ;
      END
   END n_4867

   PIN n_4868
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 20.05 0 20.15 0.51 ;
      END
   END n_4868

   PIN n_4933
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 67.65 0 67.75 0.51 ;
      END
   END n_4933

   PIN n_5261
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 0 86.95 0.51 87.05 ;
      END
   END n_5261

   PIN n_5296
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 0 63.95 0.51 64.05 ;
      END
   END n_5296

   PIN n_65597
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 15.35 280 15.45 ;
      END
   END n_65597

   PIN n_65740
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 52.15 280 52.25 ;
      END
   END n_65740

   PIN n_65860
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 63.95 280 64.05 ;
      END
   END n_65860

   PIN n_6598
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 197.05 0 197.15 0.51 ;
      END
   END n_6598

   PIN n_66080
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.745 13.3 280 13.5 ;
      END
   END n_66080

   PIN n_66260
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 75.95 280 76.05 ;
      END
   END n_66260

   PIN n_6675
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 164.05 0 164.15 0.51 ;
      END
   END n_6675

   PIN n_7855
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 163.85 0 163.95 0.51 ;
      END
   END n_7855

   PIN n_8357
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 159.85 0 159.95 0.51 ;
      END
   END n_8357

   PIN n_8586
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 158.65 0 158.75 0.51 ;
      END
   END n_8586

   PIN n_8587
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 156.45 0 156.55 0.51 ;
      END
   END n_8587

   PIN n_8743
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.25 0 115.35 0.51 ;
      END
   END n_8743

   PIN n_8902
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 131.05 0 131.15 0.51 ;
      END
   END n_8902

   PIN n_91003
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 111.35 280 111.45 ;
      END
   END n_91003

   PIN n_91051
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 279.745 11.1 280 11.3 ;
      END
   END n_91051

   PIN n_91073
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 270.65 0 270.75 0.51 ;
      END
   END n_91073

   PIN n_91091
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 100.15 280 100.25 ;
      END
   END n_91091

   PIN n_91165
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 12.95 280 13.05 ;
      END
   END n_91165

   PIN n_91268
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 272.25 0 272.35 0.51 ;
      END
   END n_91268

   PIN n_91345
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 15.15 280 15.25 ;
      END
   END n_91345

   PIN n_91373
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 274.65 0 274.75 0.51 ;
      END
   END n_91373

   PIN n_91534
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 87.75 280 87.85 ;
      END
   END n_91534

   PIN n_91579
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 12.75 280 12.85 ;
      END
   END n_91579

   PIN n_92127
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 111.95 280 112.05 ;
      END
   END n_92127

   PIN n_92142
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 111.75 280 111.85 ;
      END
   END n_92142

   PIN n_92144
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 124.15 280 124.25 ;
      END
   END n_92144

   PIN n_92271
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 88.15 280 88.25 ;
      END
   END n_92271

   PIN n_92319
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 14.95 280 15.05 ;
      END
   END n_92319

   PIN n_92482
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 111.55 280 111.65 ;
      END
   END n_92482

   PIN n_934
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 203.45 0 203.55 0.51 ;
      END
   END n_934

   PIN n_935
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 106.65 0 106.75 0.51 ;
      END
   END n_935

   PIN n_9426
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 115.05 0 115.15 0.51 ;
      END
   END n_9426

   PIN n_9428
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 155.45 0 155.55 0.51 ;
      END
   END n_9428

   PIN n_9499
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.25 0 116.35 0.51 ;
      END
   END n_9499

   PIN n_95152
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 147.55 280 147.65 ;
      END
   END n_95152

   PIN n_95239
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 135.75 280 135.85 ;
      END
   END n_95239

   PIN n_95318
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 135.55 280 135.65 ;
      END
   END n_95318

   PIN n_95323
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 14.75 280 14.85 ;
      END
   END n_95323

   PIN n_95363
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 11.95 280 12.05 ;
      END
   END n_95363

   PIN n_95397
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 14.55 280 14.65 ;
      END
   END n_95397

   PIN n_95412
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 14.35 280 14.45 ;
      END
   END n_95412

   PIN n_95416
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 14.15 280 14.25 ;
      END
   END n_95416

   PIN n_95587
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 13.95 280 14.05 ;
      END
   END n_95587

   PIN n_95604
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.745 11.5 280 11.7 ;
      END
   END n_95604

   PIN n_95698
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 147.75 280 147.85 ;
      END
   END n_95698

   PIN n_95810
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 147.95 280 148.05 ;
      END
   END n_95810

   PIN n_96003
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 159.95 280 160.05 ;
      END
   END n_96003

   PIN n_96004
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 12.55 280 12.65 ;
      END
   END n_96004

   PIN n_96232
      DIRECTION INPUT ;
      PORT 
         LAYER metal3 ;
             RECT 279.49 12.35 280 12.45 ;
      END
   END n_96232

   PIN n_96447
      DIRECTION INPUT ;
      PORT 
         LAYER metal5 ;
             RECT 279.49 11.55 280 11.65 ;
      END
   END n_96447

   PIN n_9741
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 116.05 0 116.15 0.51 ;
      END
   END n_9741

   PIN n_9764
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 140.05 0 140.15 0.51 ;
      END
   END n_9764

   PIN u0_IP_64__1294
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 212.65 0 212.75 0.51 ;
      END
   END u0_IP_64__1294

   PIN u0_R0_10_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 231.85 0 231.95 0.51 ;
      END
   END u0_R0_10_

   PIN u0_R0_20_
      DIRECTION INPUT ;
      PORT 
         LAYER metal4 ;
             RECT 206.85 0 206.95 0.51 ;
      END
   END u0_R0_20_

   PIN u0_R0_24_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 144.45 0 144.55 0.51 ;
      END
   END u0_R0_24_

   PIN u0_R0_26_
      DIRECTION INPUT ;
      PORT 
         LAYER metal2 ;
             RECT 193.25 0 193.35 0.51 ;
      END
   END u0_R0_26_

   OBS
      LAYER via4 ;
         RECT 0 0 280 296.81 ;
      LAYER via3 ;
         RECT 0 0 280 296.81 ;
      LAYER via2 ;
         RECT 0 0 280 296.81 ;
      LAYER via1 ;
         RECT 0 0 280 296.81 ;
      LAYER metal5 ;
         RECT 0 0 280 296.81 ;
      LAYER metal4 ;
         RECT 0 0 280 296.81 ;
      LAYER metal3 ;
         RECT 0 0 280 296.81 ;
      LAYER metal2 ;
         RECT 0 0 280 296.81 ;
      LAYER metal1 ;
         RECT 0 0 280 296.81 ;
   END
END h0

MACRO ms00f80
   CLASS CORE ;
   FOREIGN ms00f80 ;
   ORIGIN 0 0 ;
   SIZE 1.6 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN ck
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END ck

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.05 0.5 1.15 1.5 ;
      END
   END d

END ms00f80

MACRO in01f01
   CLASS CORE ;
   FOREIGN in01f01 ;
   ORIGIN 0 0 ;
   SIZE 0.4 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

END in01f01

MACRO na02f01
   CLASS CORE ;
   FOREIGN na02f01 ;
   ORIGIN 0 0 ;
   SIZE 0.8 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

END na02f01

MACRO no02f01
   CLASS CORE ;
   FOREIGN no02f01 ;
   ORIGIN 0 0 ;
   SIZE 0.8 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.45 0.5 0.55 1.5 ;
      END
   END b

END no02f01

MACRO oa12f01
   CLASS CORE ;
   FOREIGN oa12f01 ;
   ORIGIN 0 0 ;
   SIZE 1.2 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

END oa12f01

MACRO na04m01
   CLASS CORE ;
   FOREIGN na04m01 ;
   ORIGIN 0 0 ;
   SIZE 1.6 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

END na04m01

MACRO ao12f01
   CLASS CORE ;
   FOREIGN ao12f01 ;
   ORIGIN 0 0 ;
   SIZE 1.2 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

END ao12f01

MACRO na03f01
   CLASS CORE ;
   FOREIGN na03f01 ;
   ORIGIN 0 0 ;
   SIZE 1.2 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

END na03f01

MACRO ao22s01
   CLASS CORE ;
   FOREIGN ao22s01 ;
   ORIGIN 0 0 ;
   SIZE 1.6 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

END ao22s01

MACRO oa22f01
   CLASS CORE ;
   FOREIGN oa22f01 ;
   ORIGIN 0 0 ;
   SIZE 1.6 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal2 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

END oa22f01

MACRO no03m01
   CLASS CORE ;
   FOREIGN no03m01 ;
   ORIGIN 0 0 ;
   SIZE 1.2 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

END no03m01

MACRO no04s01
   CLASS CORE ;
   FOREIGN no04s01 ;
   ORIGIN 0 0 ;
   SIZE 1.6 BY 2 ;
   SYMMETRY X Y R90 ;
   SITE core ;
   PIN o
      DIRECTION OUTPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.05 0.5 0.15 1.5 ;
      END
   END o

   PIN a
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.25 0.5 0.35 1.5 ;
      END
   END a

   PIN b
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.65 0.5 0.75 1.5 ;
      END
   END b

   PIN c
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 0.85 0.5 0.95 1.5 ;
      END
   END c

   PIN d
      DIRECTION INPUT ;
      PORT 
         LAYER metal1 ;
             RECT 1.25 0.5 1.35 1.5 ;
      END
   END d

END no04s01

END LIBRARY
